/******************************************************************************

    File Name:  pwm_gen.v
      Version:  4.0
         Date:  July 14th, 2009
  Description:  PWM Generation Module
  
  
  SVN Revision Information:
  SVN $Revision: 10769 $
  SVN $Date: 2009-11-05 15:38:11 -0800 (Thu, 05 Nov 2009) $  
  
  

 COPYRIGHT 2009 BY ACTEL 
 THE INFORMATION CONTAINED IN THIS DOCUMENT IS SUBJECT TO LICENSING RESTRICTIONS 
 FROM ACTEL CORP.  IF YOU ARE NOT IN POSSESSION OF WRITTEN AUTHORIZATION FROM 
 ACTEL FOR USE OF THIS FILE, THEN THE FILE SHOULD BE IMMEDIATELY DESTROYED AND 
 NO BACK-UP OF THE FILE SHOULD BE MADE. 
 
FUNCTIONAL DESCRIPTION: 
Refer to the CorePWM Handbook.
******************************************************************************/
`timescale 1ns/1ns
module
pwm_gen
#
(
parameter
PWM_NUM
=
8
,
parameter
APB_DWIDTH
=
8
,
parameter
DAC_MODE
=
0
)
(
input
PRESETN,
input
PCLK,
output
[
PWM_NUM
:
1
]
PWM,
input
[
APB_DWIDTH
-
1
:
0
]
period_cnt,
input
[
PWM_NUM
:
1
]
pwm_enable_reg,
input
[
PWM_NUM
*
APB_DWIDTH
:
1
]
pwm_posedge_reg,
input
[
PWM_NUM
*
APB_DWIDTH
:
1
]
pwm_negedge_reg,
input
sync_pulse
)
;
reg
[
PWM_NUM
:
1
]
CPWMO
;
reg
[
PWM_NUM
*
(
APB_DWIDTH
+
1
)
:
1
]
CPWMOl1
;
assign
PWM
[
PWM_NUM
:
1
]
=
CPWMO
[
PWM_NUM
:
1
]
;
genvar
CPWMIl1
;
generate
for
(
CPWMIl1
=
1
;
CPWMIl1
<=
PWM_NUM
;
CPWMIl1
=
CPWMIl1
+
1
)
begin
:
CPWMll1
if
(
DAC_MODE
[
CPWMIl1
-
1
]
==
0
)
begin
always
@
(
negedge
PRESETN
or
posedge
PCLK
)
begin
if
(
!
PRESETN
)
begin
CPWMO
[
CPWMIl1
]
<=
1
'b
0
;
end
else
begin
if
(
pwm_enable_reg
[
CPWMIl1
]
==
1
'b
0
)
begin
CPWMO
[
CPWMIl1
]
<=
1
'b
0
;
end
else
if
(
(
pwm_enable_reg
[
CPWMIl1
]
==
1
'b
1
)
&&
(
sync_pulse
==
1
'b
1
)
)
begin
if
(
(
pwm_posedge_reg
[
CPWMIl1
*
APB_DWIDTH
:
(
CPWMIl1
-
1
)
*
APB_DWIDTH
+
1
]
==
pwm_negedge_reg
[
CPWMIl1
*
APB_DWIDTH
:
(
CPWMIl1
-
1
)
*
APB_DWIDTH
+
1
]
)
&&
(
(
pwm_posedge_reg
[
CPWMIl1
*
APB_DWIDTH
:
(
CPWMIl1
-
1
)
*
APB_DWIDTH
+
1
]
)
==
period_cnt
)
)
begin
CPWMO
[
CPWMIl1
]
<=
~
CPWMO
[
CPWMIl1
]
;
end
else
if
(
(
pwm_enable_reg
[
CPWMIl1
]
==
1
'b
1
)
&&
(
sync_pulse
==
1
'b
1
)
&&
(
pwm_posedge_reg
[
CPWMIl1
*
APB_DWIDTH
:
(
CPWMIl1
-
1
)
*
APB_DWIDTH
+
1
]
)
==
period_cnt
)
begin
CPWMO
[
CPWMIl1
]
<=
1
'b
1
;
end
else
if
(
(
pwm_enable_reg
[
CPWMIl1
]
==
1
'b
1
)
&&
(
sync_pulse
==
1
'b
1
)
&&
(
pwm_negedge_reg
[
CPWMIl1
*
APB_DWIDTH
:
(
CPWMIl1
-
1
)
*
APB_DWIDTH
+
1
]
)
==
period_cnt
)
begin
CPWMO
[
CPWMIl1
]
<=
1
'b
0
;
end
end
end
end
end
else
begin
always
@
(
negedge
PRESETN
or
posedge
PCLK
)
begin
if
(
!
PRESETN
)
begin
CPWMOl1
[
CPWMIl1
*
(
APB_DWIDTH
+
1
)
:
(
CPWMIl1
-
1
)
*
(
APB_DWIDTH
+
1
)
+
1
]
<=
0
;
CPWMO
[
CPWMIl1
]
<=
1
'b
0
;
end
else
begin
if
(
pwm_enable_reg
[
CPWMIl1
]
==
1
'b
0
)
begin
CPWMO
[
CPWMIl1
]
<=
1
'b
0
;
end
else
if
(
pwm_enable_reg
[
CPWMIl1
]
==
1
'b
1
)
begin
CPWMOl1
[
CPWMIl1
*
(
APB_DWIDTH
+
1
)
:
(
CPWMIl1
-
1
)
*
(
APB_DWIDTH
+
1
)
+
1
]
<=
CPWMOl1
[
(
CPWMIl1
*
(
APB_DWIDTH
+
1
)
)
-
1
:
(
CPWMIl1
-
1
)
*
(
APB_DWIDTH
+
1
)
+
1
]
+
pwm_negedge_reg
[
CPWMIl1
*
APB_DWIDTH
:
(
CPWMIl1
-
1
)
*
APB_DWIDTH
+
1
]
;
CPWMO
[
CPWMIl1
]
<=
CPWMOl1
[
CPWMIl1
*
(
APB_DWIDTH
+
1
)
]
;
end
end
end
end
end
endgenerate
endmodule
