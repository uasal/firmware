// Actel Corporation Proprietary and Confidential
// Copyright 2013 Actel Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE ACTEL LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
// SVN Revision Information:
// SVN $Revision: 23120 $
// SVN $Date: 2014-07-17 15:26:23 +0100 (Thu, 17 Jul 2014) $
`timescale 1ns/1ps
module
CAHBLTOI1I
#
(
parameter
SYNC_RESET
=
0
)
(
input
HCLK,
input
HRESETN,
input
CAHBLTII1I,
input
CAHBLTI0OI,
output
reg
CAHBLTlI1I,
output
reg
[
31
:
0
]
CAHBLTlIOI,
output
reg
[
2
:
0
]
CAHBLTIlOI,
output
wire
CAHBLTllOI,
output
reg
CAHBLTO0OI,
output
reg
[
31
:
0
]
CAHBLTOl1I,
output
wire
CAHBLTIl1I,
output
reg
CAHBLTOlOI,
input
[
3
:
0
]
CAHBLTOI0,
input
[
3
:
0
]
CAHBLTll1I,
input
[
3
:
0
]
CAHBLTO01I,
output
reg
[
3
:
0
]
CAHBLTI01I,
output
reg
[
3
:
0
]
CAHBLTl01I,
output
reg
[
3
:
0
]
CAHBLTO11I,
input
[
31
:
0
]
CAHBLTI11I,
input
CAHBLTlI0,
input
[
2
:
0
]
CAHBLTl11I,
input
CAHBLTOOOl,
input
CAHBLTIOOl,
input
[
31
:
0
]
CAHBLTlOOl,
input
CAHBLTOl0,
input
[
2
:
0
]
CAHBLTOIOl,
input
CAHBLTIIOl,
input
CAHBLTlIOl,
input
[
31
:
0
]
CAHBLTOlOl,
input
CAHBLTIl0,
input
[
2
:
0
]
CAHBLTIlOl,
input
CAHBLTllOl,
input
CAHBLTO0Ol,
input
[
31
:
0
]
CAHBLTI0Ol,
input
CAHBLTll0,
input
[
2
:
0
]
CAHBLTl0Ol,
input
CAHBLTO1Ol,
input
CAHBLTI1Ol,
input
[
31
:
0
]
HWDATA_M0,
input
[
31
:
0
]
HWDATA_M1,
input
[
31
:
0
]
HWDATA_M2,
input
[
31
:
0
]
HWDATA_M3
)
;
localparam
CAHBLTl1Ol
=
1
'b
0
;
localparam
CAHBLTOOOI
=
4
'b
0000
;
wire
[
3
:
0
]
CAHBLTOOIl
;
reg
[
3
:
0
]
CAHBLTIOIl
;
reg
CAHBLTlOIl
;
wire
CAHBLTOIIl
;
reg
CAHBLTIIIl
;
wire
CAHBLTOO0
;
wire
CAHBLTIO0
;
assign
CAHBLTOO0
=
(
SYNC_RESET
==
1
)
?
1
'b
1
:
HRESETN
;
assign
CAHBLTIO0
=
(
SYNC_RESET
==
1
)
?
HRESETN
:
1
'b
1
;
always
@
(
posedge
HCLK
or
negedge
CAHBLTOO0
)
begin
if
(
(
!
CAHBLTOO0
)
||
(
!
CAHBLTIO0
)
)
CAHBLTIOIl
<=
CAHBLTOOOI
;
else
if
(
CAHBLTIl1I
)
CAHBLTIOIl
<=
CAHBLTOOIl
;
end
CAHBLTlO0
#
(
.SYNC_RESET
(
SYNC_RESET
)
)
CAHBLTlIIl
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.CAHBLTOI0
(
CAHBLTOI0
)
,
.CAHBLTII0
(
CAHBLTIl1I
)
,
.CAHBLTlI0
(
CAHBLTlI0
)
,
.CAHBLTOl0
(
CAHBLTOl0
)
,
.CAHBLTIl0
(
CAHBLTIl0
)
,
.CAHBLTll0
(
CAHBLTll0
)
,
.CAHBLTO00
(
CAHBLTOOIl
)
)
;
always
@
(
*
)
begin
casez
(
CAHBLTOOIl
)
4
'b
???1
:
begin
CAHBLTlI1I
=
1
'b
1
;
CAHBLTIIIl
=
CAHBLTOOOl
;
CAHBLTIlOI
=
CAHBLTl11I
;
CAHBLTO0OI
=
CAHBLTIOOl
;
CAHBLTlIOI
=
CAHBLTI11I
;
CAHBLTOlOI
=
CAHBLTlI0
;
CAHBLTlOIl
=
CAHBLTO01I
[
0
]
;
end
4
'b
??1?
:
begin
CAHBLTlI1I
=
1
'b
1
;
CAHBLTIIIl
=
CAHBLTIIOl
;
CAHBLTIlOI
=
CAHBLTOIOl
;
CAHBLTO0OI
=
CAHBLTlIOl
;
CAHBLTlIOI
=
CAHBLTlOOl
;
CAHBLTOlOI
=
CAHBLTOl0
;
CAHBLTlOIl
=
CAHBLTO01I
[
1
]
;
end
4
'b
?1??
:
begin
CAHBLTlI1I
=
1
'b
1
;
CAHBLTIIIl
=
CAHBLTllOl
;
CAHBLTIlOI
=
CAHBLTIlOl
;
CAHBLTO0OI
=
CAHBLTO0Ol
;
CAHBLTlIOI
=
CAHBLTOlOl
;
CAHBLTOlOI
=
CAHBLTIl0
;
CAHBLTlOIl
=
CAHBLTO01I
[
2
]
;
end
4
'b
1???
:
begin
CAHBLTlI1I
=
1
'b
1
;
CAHBLTIIIl
=
CAHBLTO1Ol
;
CAHBLTIlOI
=
CAHBLTl0Ol
;
CAHBLTO0OI
=
CAHBLTI1Ol
;
CAHBLTlIOI
=
CAHBLTI0Ol
;
CAHBLTOlOI
=
CAHBLTll0
;
CAHBLTlOIl
=
CAHBLTO01I
[
3
]
;
end
default
:
begin
CAHBLTlI1I
=
1
'b
0
;
CAHBLTIIIl
=
CAHBLTl1Ol
;
CAHBLTIlOI
=
2
'b
00
;
CAHBLTO0OI
=
1
'b
0
;
CAHBLTlIOI
=
32
'h
0
;
CAHBLTOlOI
=
1
'b
0
;
CAHBLTlOIl
=
1
'b
1
;
end
endcase
end
assign
CAHBLTOIIl
=
|
(
CAHBLTOOIl
&
CAHBLTll1I
)
;
assign
CAHBLTllOI
=
CAHBLTIIIl
&&
(
CAHBLTlOIl
||
CAHBLTOIIl
)
;
assign
CAHBLTIl1I
=
CAHBLTII1I
;
always
@
(
*
)
begin
casez
(
CAHBLTIOIl
)
4
'b
???1
:
begin
CAHBLTOl1I
=
HWDATA_M0
;
end
4
'b
??1?
:
begin
CAHBLTOl1I
=
HWDATA_M1
;
end
4
'b
?1??
:
begin
CAHBLTOl1I
=
HWDATA_M2
;
end
4
'b
1???
:
begin
CAHBLTOl1I
=
HWDATA_M3
;
end
default
:
begin
CAHBLTOl1I
=
32
'h
0
;
end
endcase
end
always
@
(
*
)
begin
CAHBLTO11I
=
2
'b
00
;
casez
(
CAHBLTIOIl
)
4
'b
???1
:
begin
CAHBLTO11I
[
0
]
=
CAHBLTI0OI
;
end
4
'b
??1?
:
begin
CAHBLTO11I
[
1
]
=
CAHBLTI0OI
;
end
4
'b
?1??
:
begin
CAHBLTO11I
[
2
]
=
CAHBLTI0OI
;
end
4
'b
1???
:
begin
CAHBLTO11I
[
3
]
=
CAHBLTI0OI
;
end
default
:
begin
CAHBLTO11I
=
2
'b
00
;
end
endcase
end
always
@
(
*
)
begin
if
(
CAHBLTOI0
[
0
]
&&
!
CAHBLTOOIl
[
0
]
)
CAHBLTI01I
[
0
]
=
1
'b
0
;
else
if
(
CAHBLTOI0
[
0
]
&&
CAHBLTOOIl
[
0
]
)
CAHBLTI01I
[
0
]
=
CAHBLTII1I
;
else
CAHBLTI01I
[
0
]
=
1
'b
1
;
end
always
@
(
*
)
begin
if
(
CAHBLTOI0
[
1
]
&&
!
CAHBLTOOIl
[
1
]
)
CAHBLTI01I
[
1
]
=
1
'b
0
;
else
if
(
CAHBLTOI0
[
1
]
&&
CAHBLTOOIl
[
1
]
)
CAHBLTI01I
[
1
]
=
CAHBLTII1I
;
else
CAHBLTI01I
[
1
]
=
1
'b
1
;
end
always
@
(
*
)
begin
if
(
CAHBLTOI0
[
2
]
&&
!
CAHBLTOOIl
[
2
]
)
CAHBLTI01I
[
2
]
=
1
'b
0
;
else
if
(
CAHBLTOI0
[
2
]
&&
CAHBLTOOIl
[
2
]
)
CAHBLTI01I
[
2
]
=
CAHBLTII1I
;
else
CAHBLTI01I
[
2
]
=
1
'b
1
;
end
always
@
(
*
)
begin
if
(
CAHBLTOI0
[
3
]
&&
!
CAHBLTOOIl
[
3
]
)
CAHBLTI01I
[
3
]
=
1
'b
0
;
else
if
(
CAHBLTOI0
[
3
]
&&
CAHBLTOOIl
[
3
]
)
CAHBLTI01I
[
3
]
=
CAHBLTII1I
;
else
CAHBLTI01I
[
3
]
=
1
'b
1
;
end
always
@
(
*
)
begin
if
(
CAHBLTll1I
[
0
]
&&
!
CAHBLTIOIl
[
0
]
)
CAHBLTl01I
[
0
]
=
1
'b
0
;
else
if
(
CAHBLTll1I
[
0
]
&&
CAHBLTIOIl
[
0
]
)
CAHBLTl01I
[
0
]
=
CAHBLTII1I
;
else
CAHBLTl01I
[
0
]
=
1
'b
1
;
end
always
@
(
*
)
begin
if
(
CAHBLTll1I
[
1
]
&&
!
CAHBLTIOIl
[
1
]
)
CAHBLTl01I
[
1
]
=
1
'b
0
;
else
if
(
CAHBLTll1I
[
1
]
&&
CAHBLTIOIl
[
1
]
)
CAHBLTl01I
[
1
]
=
CAHBLTII1I
;
else
CAHBLTl01I
[
1
]
=
1
'b
1
;
end
always
@
(
*
)
begin
if
(
CAHBLTll1I
[
2
]
&&
!
CAHBLTIOIl
[
2
]
)
CAHBLTl01I
[
2
]
=
1
'b
0
;
else
if
(
CAHBLTll1I
[
2
]
&&
CAHBLTIOIl
[
2
]
)
CAHBLTl01I
[
2
]
=
CAHBLTII1I
;
else
CAHBLTl01I
[
2
]
=
1
'b
1
;
end
always
@
(
*
)
begin
if
(
CAHBLTll1I
[
3
]
&&
!
CAHBLTIOIl
[
3
]
)
CAHBLTl01I
[
3
]
=
1
'b
0
;
else
if
(
CAHBLTll1I
[
3
]
&&
CAHBLTIOIl
[
3
]
)
CAHBLTl01I
[
3
]
=
CAHBLTII1I
;
else
CAHBLTl01I
[
3
]
=
1
'b
1
;
end
endmodule
