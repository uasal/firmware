-- megafunction wizard: %Altera Unique Chip ID v14.1%
-- GENERATION: XML
-- Serial.vhd

-- Generated using ACDS version 14.1 186 at 2015.11.13.16:00:02

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Serial is
	port (
		clkin      : in  std_logic                     := '0'; --  clkin.clk
		reset      : in  std_logic                     := '0'; --  reset.reset
		data_valid : out std_logic;                            -- output.valid
		chip_id    : out std_logic_vector(63 downto 0)         --       .data
	);
end entity Serial;

architecture rtl of Serial is
	component altchip_id is
		generic (
			DEVICE_FAMILY : string                        := "";
			ID_VALUE      : std_logic_vector(63 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111";
			ID_VALUE_STR  : string                        := "ffffffffffffffff"
		);
		port (
			clkin      : in  std_logic                     := 'X'; -- clk
			reset      : in  std_logic                     := 'X'; -- reset
			data_valid : out std_logic;                            -- valid
			chip_id    : out std_logic_vector(63 downto 0)         -- data
		);
	end component altchip_id;

begin

	serial_inst : component altchip_id
		generic map (
			DEVICE_FAMILY => "MAX 10",
			ID_VALUE      => "1111111111111111111111111111111111111111111111111111111111111111",
			ID_VALUE_STR  => "ffffffffffffffff"
		)
		port map (
			clkin      => clkin,      --  clkin.clk
			reset      => reset,      --  reset.reset
			data_valid => data_valid, -- output.valid
			chip_id    => chip_id     --       .data
		);

end architecture rtl; -- of Serial
-- Retrieval info: <?xml version="1.0"?>
--<!--
--	Generated by Altera MegaWizard Launcher Utility version 1.0
--	************************************************************
--	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--	************************************************************
--	Copyright (C) 1991-2015 Altera Corporation
--	Any megafunction design, and related net list (encrypted or decrypted),
--	support information, device programming or simulation file, and any other
--	associated documentation or information provided by Altera or a partner
--	under Altera's Megafunction Partnership Program may be used only to
--	program PLD devices (but not masked PLD devices) from Altera.  Any other
--	use of such megafunction design, net list, support information, device
--	programming or simulation file, or any other related documentation or
--	information is prohibited for any other purpose, including, but not
--	limited to modification, reverse engineering, de-compiling, or use with
--	any other silicon devices, unless such use is explicitly licensed under
--	a separate agreement with Altera or a megafunction partner.  Title to
--	the intellectual property, including patents, copyrights, trademarks,
--	trade secrets, or maskworks, embodied in any such megafunction design,
--	net list, support information, device programming or simulation file, or
--	any other related documentation or information provided by Altera or a
--	megafunction partner, remains with Altera, the megafunction partner, or
--	their respective licensors.  No other licenses, including any licenses
--	needed under any third party's intellectual property, are provided herein.
---->
-- Retrieval info: <instance entity-name="altchip_id" version="14.1" >
-- Retrieval info: 	<generic name="DEVICE_FAMILY" value="MAX 10" />
-- Retrieval info: 	<generic name="ID_VALUE" value="18446744073709551615" />
-- Retrieval info: </instance>
-- IPFS_FILES : Serial.vho
-- RELATED_FILES: Serial.vhd, altchip_id.v
