// Actel Corporation Proprietary and Confidential
// Copyright 2010 Actel Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE ACTEL LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
// SVN Revision Information:
// SVN $Revision: 23120 $
// SVN $Date: 2014-07-17 15:26:23 +0100 (Thu, 17 Jul 2014) $
`timescale 1ns/1ps
module
CAHBLTO
#
(
parameter
[
2
:
0
]
MEMSPACE
=
0
,
parameter
[
0
:
0
]
HADDR_SHG_CFG
=
1
,
parameter
[
15
:
0
]
CAHBLTI
=
0
,
parameter
[
16
:
0
]
CAHBLTl
=
(
2
**
17
)
-
1
)
(
input
[
31
:
0
]
CAHBLTOI,
input
CAHBLTII,
output
wire
[
16
:
0
]
CAHBLTlI,
output
wire
[
31
:
0
]
CAHBLTOl,
output
wire
CAHBLTIl
)
;
localparam
CAHBLTll
=
(
MEMSPACE
==
1
)
?
31
:
(
MEMSPACE
==
2
)
?
27
:
(
MEMSPACE
==
3
)
?
23
:
(
MEMSPACE
==
4
)
?
19
:
(
MEMSPACE
==
5
)
?
15
:
(
MEMSPACE
==
6
)
?
11
:
31
;
localparam
CAHBLTO0
=
16
'b
0000000000000001
;
localparam
CAHBLTI0
=
16
'b
0000000000000010
;
localparam
CAHBLTl0
=
16
'b
0000000000000100
;
localparam
CAHBLTO1
=
16
'b
0000000000001000
;
localparam
CAHBLTI1
=
16
'b
0000000000010000
;
localparam
CAHBLTl1
=
16
'b
0000000000100000
;
localparam
CAHBLTOOI
=
16
'b
0000000001000000
;
localparam
CAHBLTIOI
=
16
'b
0000000010000000
;
localparam
CAHBLTlOI
=
16
'b
0000000100000000
;
localparam
CAHBLTOII
=
16
'b
0000001000000000
;
localparam
CAHBLTIII
=
16
'b
0000010000000000
;
localparam
CAHBLTlII
=
16
'b
0000100000000000
;
localparam
CAHBLTOlI
=
16
'b
0001000000000000
;
localparam
CAHBLTIlI
=
16
'b
0010000000000000
;
localparam
CAHBLTllI
=
16
'b
0100000000000000
;
localparam
CAHBLTO0I
=
16
'b
1000000000000000
;
localparam
CAHBLTI0I
=
16
'b
0000000000000000
;
reg
[
15
:
0
]
CAHBLTl0I
;
reg
[
15
:
0
]
CAHBLTO1I
;
reg
CAHBLTI1I
;
reg
[
31
:
0
]
CAHBLTl1I
;
wire
[
16
:
0
]
CAHBLTOOl
;
wire
[
3
:
0
]
CAHBLTIOl
;
wire
CAHBLTlOl
;
wire
CAHBLTOIl
;
generate
begin
:
CAHBLTIIl
if
(
MEMSPACE
==
0
)
begin
:
CAHBLTlIl
assign
CAHBLTlOl
=
(
CAHBLTOI
[
31
]
==
1
'b
1
)
;
assign
CAHBLTOIl
=
(
CAHBLTOI
[
30
:
20
]
==
11
'h
000
)
;
assign
CAHBLTIOl
=
CAHBLTOI
[
19
:
16
]
;
always
@
(
*
)
begin
CAHBLTl1I
[
31
:
0
]
=
CAHBLTOI
[
31
:
0
]
;
CAHBLTl0I
[
15
:
0
]
=
CAHBLTI0I
;
if
(
CAHBLTlOl
)
begin
CAHBLTI1I
=
1
'b
1
;
if
(
HADDR_SHG_CFG
==
0
)
begin
CAHBLTl1I
[
31
]
=
1
'b
0
;
end
else
begin
CAHBLTl1I
[
31
]
=
1
'b
1
;
end
end
else
if
(
CAHBLTOIl
)
begin
case
(
CAHBLTIOl
)
4
'h
0
:
begin
if
(
CAHBLTII
==
1
'b
0
)
begin
CAHBLTl0I
[
15
:
0
]
=
CAHBLTO0
;
end
else
begin
CAHBLTl1I
[
16
]
=
1
'b
1
;
CAHBLTl0I
[
15
:
0
]
=
CAHBLTI0
;
end
end
4
'h
1
:
begin
if
(
CAHBLTII
==
1
'b
0
)
begin
CAHBLTl0I
[
15
:
0
]
=
CAHBLTI0
;
end
else
begin
CAHBLTl1I
[
16
]
=
1
'b
0
;
CAHBLTl0I
[
15
:
0
]
=
CAHBLTO0
;
end
end
4
'h
2
:
CAHBLTl0I
[
15
:
0
]
=
CAHBLTl0
;
4
'h
3
:
CAHBLTl0I
[
15
:
0
]
=
CAHBLTO1
;
4
'h
4
:
CAHBLTl0I
[
15
:
0
]
=
CAHBLTI1
;
4
'h
5
:
CAHBLTl0I
[
15
:
0
]
=
CAHBLTl1
;
4
'h
6
:
CAHBLTl0I
[
15
:
0
]
=
CAHBLTOOI
;
4
'h
7
:
CAHBLTl0I
[
15
:
0
]
=
CAHBLTIOI
;
4
'h
8
:
CAHBLTl0I
[
15
:
0
]
=
CAHBLTlOI
;
4
'h
9
:
CAHBLTl0I
[
15
:
0
]
=
CAHBLTOII
;
4
'h
A
:
CAHBLTl0I
[
15
:
0
]
=
CAHBLTIII
;
4
'h
B
:
CAHBLTl0I
[
15
:
0
]
=
CAHBLTlII
;
4
'h
C
:
CAHBLTl0I
[
15
:
0
]
=
CAHBLTOlI
;
4
'h
D
:
CAHBLTl0I
[
15
:
0
]
=
CAHBLTIlI
;
4
'h
E
:
CAHBLTl0I
[
15
:
0
]
=
CAHBLTllI
;
4
'h
F
:
CAHBLTl0I
[
15
:
0
]
=
CAHBLTO0I
;
endcase
end
CAHBLTO1I
=
CAHBLTl0I
;
CAHBLTI1I
=
CAHBLTlOl
;
end
assign
CAHBLTIl
=
CAHBLTlOl
==
1
'b
0
&
CAHBLTOIl
==
1
'b
0
;
end
else
begin
:
CAHBLTOll
assign
CAHBLTlOl
=
1
'b
0
;
assign
CAHBLTOIl
=
1
'b
0
;
assign
CAHBLTIOl
=
CAHBLTOI
[
CAHBLTll
:
CAHBLTll
-
3
]
;
always
@
(
*
)
begin
CAHBLTl1I
[
31
:
0
]
=
CAHBLTOI
[
31
:
0
]
;
case
(
CAHBLTIOl
)
4
'h
0
:
begin
if
(
CAHBLTII
==
1
'b
0
)
CAHBLTl0I
[
15
:
0
]
=
CAHBLTO0
;
else
begin
CAHBLTl1I
[
CAHBLTll
-
3
]
=
1
'b
1
;
CAHBLTl0I
[
15
:
0
]
=
CAHBLTI0
;
end
end
4
'h
1
:
begin
if
(
CAHBLTII
==
1
'b
0
)
CAHBLTl0I
[
15
:
0
]
=
CAHBLTI0
;
else
begin
CAHBLTl1I
[
CAHBLTll
-
3
]
=
1
'b
0
;
CAHBLTl0I
[
15
:
0
]
=
CAHBLTO0
;
end
end
4
'h
2
:
CAHBLTl0I
[
15
:
0
]
=
CAHBLTl0
;
4
'h
3
:
CAHBLTl0I
[
15
:
0
]
=
CAHBLTO1
;
4
'h
4
:
CAHBLTl0I
[
15
:
0
]
=
CAHBLTI1
;
4
'h
5
:
CAHBLTl0I
[
15
:
0
]
=
CAHBLTl1
;
4
'h
6
:
CAHBLTl0I
[
15
:
0
]
=
CAHBLTOOI
;
4
'h
7
:
CAHBLTl0I
[
15
:
0
]
=
CAHBLTIOI
;
4
'h
8
:
CAHBLTl0I
[
15
:
0
]
=
CAHBLTlOI
;
4
'h
9
:
CAHBLTl0I
[
15
:
0
]
=
CAHBLTOII
;
4
'h
A
:
CAHBLTl0I
[
15
:
0
]
=
CAHBLTIII
;
4
'h
B
:
CAHBLTl0I
[
15
:
0
]
=
CAHBLTlII
;
4
'h
C
:
CAHBLTl0I
[
15
:
0
]
=
CAHBLTOlI
;
4
'h
D
:
CAHBLTl0I
[
15
:
0
]
=
CAHBLTIlI
;
4
'h
E
:
CAHBLTl0I
[
15
:
0
]
=
CAHBLTllI
;
4
'h
F
:
CAHBLTl0I
[
15
:
0
]
=
CAHBLTO0I
;
endcase
CAHBLTO1I
=
CAHBLTl0I
&
~
CAHBLTI
;
CAHBLTI1I
=
|
(
CAHBLTl0I
&
CAHBLTI
)
;
end
assign
CAHBLTIl
=
1
'b
0
;
end
assign
CAHBLTOOl
[
16
:
0
]
=
{
CAHBLTI1I
,
CAHBLTO1I
[
15
:
0
]
}
;
assign
CAHBLTOl
[
31
:
0
]
=
CAHBLTl1I
[
31
:
0
]
;
assign
CAHBLTlI
[
16
:
0
]
=
CAHBLTOOl
[
16
:
0
]
;
end
endgenerate
endmodule
