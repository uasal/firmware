//  Copyright 2011 Actel Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE ACTEL LICENSE AGREEMENT AND MUST BE APPROVED
// Revision Information:
// SVN Revision Information:
// SVN $Revision: 4805 $
`timescale 1ns/100ps
module
CHTOLSRAMII
(
HCLK
,
HRESETN
,
HSEL
,
HTRANS
,
HBURST
,
HWRITE
,
HSIZE
,
HADDR
,
HWDATA
,
HREADYIN
,
CHTOLSRAMoI
,
CHTOLSRAMOI
,
HRESP
,
HREADYOUT
,
HRDATA
,
CHTOLSRAMiI
,
CHTOLSRAMi
,
CHTOLSRAMo
,
CHTOLSRAMI
,
CHTOLSRAMl
,
BUSY
)
;
localparam
CHTOLSRAMIl
=
2
'b
00
;
localparam
CHTOLSRAMll
=
2
'b
01
;
localparam
CHTOLSRAMol
=
2
'b
10
;
parameter
AHB_DWIDTH
=
32
;
parameter
AHB_AWIDTH
=
32
;
parameter
CHTOLSRAMil
=
2
'b
00
;
parameter
CHTOLSRAMO0
=
2
'b
01
;
parameter
CHTOLSRAMI0
=
2
'b
00
;
parameter
CHTOLSRAMl0
=
2
'b
01
;
parameter
CHTOLSRAMo0
=
2
'b
11
;
parameter
CHTOLSRAMi0
=
2
'b
10
;
input
HCLK
;
input
HRESETN
;
input
HSEL
;
input
HREADYIN
;
input
[
1
:
0
]
HTRANS
;
input
[
2
:
0
]
HBURST
;
input
[
2
:
0
]
HSIZE
;
input
[
19
:
0
]
HADDR
;
input
[
AHB_DWIDTH
-
1
:
0
]
HWDATA
;
input
HWRITE
;
input
CHTOLSRAMoI
;
input
[
AHB_DWIDTH
-
1
:
0
]
CHTOLSRAMOI
;
input
BUSY
;
output
HREADYOUT
;
output
[
1
:
0
]
HRESP
;
output
[
AHB_DWIDTH
-
1
:
0
]
HRDATA
;
output
CHTOLSRAMiI
;
output
CHTOLSRAMi
;
output
[
AHB_AWIDTH
-
1
:
0
]
CHTOLSRAMo
;
output
[
2
:
0
]
CHTOLSRAMI
;
output
[
19
:
0
]
CHTOLSRAMl
;
reg
[
1
:
0
]
CHTOLSRAMO1
;
reg
[
2
:
0
]
CHTOLSRAMI1
;
reg
[
2
:
0
]
CHTOLSRAMl1
;
reg
[
19
:
0
]
CHTOLSRAMo1
;
reg
[
AHB_DWIDTH
-
1
:
0
]
CHTOLSRAMi1
;
reg
CHTOLSRAMOo
;
reg
CHTOLSRAMIo
;
reg
CHTOLSRAMlo
;
reg
[
1
:
0
]
CHTOLSRAMoo
;
reg
[
1
:
0
]
CHTOLSRAMio
;
reg
CHTOLSRAMOi
;
reg
CHTOLSRAMIi
;
reg
CHTOLSRAMli
;
reg
[
AHB_DWIDTH
-
1
:
0
]
CHTOLSRAMoi
;
reg
[
AHB_DWIDTH
-
1
:
0
]
HRDATA
;
wire
HREADYOUT
;
wire
CHTOLSRAMiI
;
wire
CHTOLSRAMii
;
wire
[
1
:
0
]
HRESP
;
wire
CHTOLSRAMi
;
wire
[
2
:
0
]
CHTOLSRAMI
;
wire
[
19
:
0
]
CHTOLSRAMl
;
assign
CHTOLSRAMii
=
HREADYIN
&
HSEL
&
(
HTRANS
==
CHTOLSRAMi0
)
;
assign
HRESP
=
CHTOLSRAMil
;
always
@
(
*
)
begin
CHTOLSRAMoi
=
HWDATA
;
end
always
@
(
posedge
HCLK
or
negedge
HRESETN
)
begin
if
(
HRESETN
==
1
'b
0
)
begin
CHTOLSRAMo1
<=
{
20
{
1
'b
0
}
}
;
CHTOLSRAMi1
<=
{
32
{
1
'b
0
}
}
;
CHTOLSRAMO1
<=
2
'b
00
;
CHTOLSRAMl1
<=
2
'b
00
;
CHTOLSRAMI1
<=
3
'b
000
;
CHTOLSRAMOo
<=
1
'b
0
;
CHTOLSRAMIo
<=
1
'b
0
;
CHTOLSRAMlo
<=
1
'b
0
;
end
else
if
(
CHTOLSRAMOi
==
1
'b
1
)
begin
CHTOLSRAMo1
<=
HADDR
;
CHTOLSRAMO1
<=
HTRANS
;
CHTOLSRAMl1
<=
HSIZE
;
CHTOLSRAMI1
<=
HBURST
;
CHTOLSRAMOo
<=
HWRITE
;
CHTOLSRAMi1
<=
CHTOLSRAMoi
;
CHTOLSRAMIo
<=
HSEL
;
CHTOLSRAMlo
<=
HREADYIN
;
end
end
always
@
(
posedge
HCLK
or
negedge
HRESETN
)
begin
if
(
HRESETN
==
1
'b
0
)
begin
CHTOLSRAMoo
<=
CHTOLSRAMIl
;
end
else
begin
CHTOLSRAMoo
<=
CHTOLSRAMio
;
end
end
always
@
(
*
)
begin
CHTOLSRAMOi
=
1
'b
0
;
CHTOLSRAMIi
=
1
'b
0
;
CHTOLSRAMio
=
CHTOLSRAMoo
;
case
(
CHTOLSRAMoo
)
CHTOLSRAMIl
:
begin
if
(
CHTOLSRAMii
==
1
'b
1
)
begin
CHTOLSRAMOi
=
1
'b
1
;
if
(
HWRITE
==
1
'b
1
)
begin
CHTOLSRAMio
=
CHTOLSRAMll
;
end
else
begin
CHTOLSRAMio
=
CHTOLSRAMol
;
end
end
end
CHTOLSRAMll
:
begin
CHTOLSRAMOi
=
1
'b
0
;
CHTOLSRAMIi
=
1
'b
1
;
if
(
CHTOLSRAMoI
==
1
'b
1
)
begin
CHTOLSRAMio
=
CHTOLSRAMIl
;
end
end
CHTOLSRAMol
:
begin
CHTOLSRAMOi
=
1
'b
0
;
CHTOLSRAMIi
=
1
'b
1
;
if
(
CHTOLSRAMoI
==
1
'b
1
)
begin
CHTOLSRAMio
=
CHTOLSRAMIl
;
end
end
default
:
begin
CHTOLSRAMio
=
CHTOLSRAMIl
;
end
endcase
end
assign
HREADYOUT
=
!
CHTOLSRAMIi
;
assign
CHTOLSRAMi
=
(
CHTOLSRAMiI
&
!
CHTOLSRAMoI
)
?
CHTOLSRAMOo
:
1
'b
0
;
assign
CHTOLSRAMo
=
HWDATA
;
assign
CHTOLSRAMl
=
(
CHTOLSRAMIi
&
!
CHTOLSRAMoI
)
?
CHTOLSRAMo1
:
CHTOLSRAMo1
;
assign
CHTOLSRAMI
=
(
CHTOLSRAMIi
&
!
CHTOLSRAMoI
)
?
CHTOLSRAMl1
:
HSIZE
;
always
@
(
posedge
HCLK
or
negedge
HRESETN
)
begin
if
(
HRESETN
==
1
'b
0
)
begin
CHTOLSRAMli
<=
1
'b
0
;
end
else
begin
CHTOLSRAMli
<=
CHTOLSRAMIi
;
end
end
assign
CHTOLSRAMiI
=
CHTOLSRAMIi
&
!
CHTOLSRAMli
&
(
CHTOLSRAMI1
==
3
'b
000
)
;
always
@
(
*
)
begin
if
(
HREADYOUT
&&
HREADYIN
)
begin
HRDATA
=
CHTOLSRAMOI
;
end
else
begin
HRDATA
=
CHTOLSRAMOI
;
end
end
endmodule
