--
--           Copyright (c) by Franks Development, LLC
--
-- This software is copyrighted by and is the sole property of Franks
-- Development, LLC. All rights, title, ownership, or other interests
-- in the software remain the property of Franks Development, LLC. This
-- software may only be used in accordance with the corresponding
-- license agreement.  Any unauthorized use, duplication, transmission,
-- distribution, or disclosure of this software is expressly forbidden.
--
-- This Copyright notice may not be removed or modified without prior
-- written consent of Franks Development, LLC.
--
-- Franks Development, LLC. reserves the right to modify this software
-- without notice.
--
-- Franks Development, LLC            support@franks-development.com
-- 500 N. Bahamas Dr. #101           http:--www.franks-development.com
-- Tucson, AZ 85710
-- USA
--
-- Permission granted for perpetual non-exclusive end-use by the University of Arizona August 1, 2020
--

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.all;
library UNISIM;
use UNISIM.vcomponents.all;

entity IOBufP3Ports is
	port (
			clk : in std_logic;
			IO  : inout std_logic;
			T : in std_logic;
			I : in std_logic;
			O : out std_logic--;
	);
end IOBufP3Ports;

architecture IOBufP3 of IOBufP3Ports is

	signal Temp1 : std_logic;
	signal Temp2 : std_logic;
	signal Temp3 : std_logic;
	
begin

	IOBUF_i : IOBUF
	port map (
		O => Temp1,
		IO => IO,
		I => I,
		T => T
	);

	process (clk)
	begin
	
		if ( (clk'event) and (clk = '1') ) then
		
			Temp2 <= Temp1; --first pipeline stage - temp2 signal
			Temp3 <= Temp2; --second pipeline stage - temp3 signal
			O <= Temp3; --third pipeline stage - O signal

		end if;

	end process; --(clock)

end IOBufP3;
