// Actel Corporation Proprietary and Confidential
// Copyright 2010 Actel Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE ACTEL LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
// SVN Revision Information:
// SVN $Revision: 23120 $
// SVN $Date: 2014-07-17 15:26:23 +0100 (Thu, 17 Jul 2014) $
`timescale 1ns/1ps
module
CAHBLTIIOI
#
(
parameter
[
2
:
0
]
MEMSPACE
=
0
,
parameter
[
0
:
0
]
HADDR_SHG_CFG
=
1
,
parameter
[
15
:
0
]
CAHBLTI
=
0
,
parameter
[
16
:
0
]
CAHBLTl
=
(
2
**
17
)
-
1
,
parameter
SYNC_RESET
=
0
)
(
input
HCLK,
input
HRESETN,
input
[
31
:
0
]
CAHBLTlIOI,
input
CAHBLTOlOI,
input
[
2
:
0
]
CAHBLTIlOI,
input
CAHBLTllOI,
input
CAHBLTO0OI,
output
reg
CAHBLTI0OI,
output
reg
[
31
:
0
]
CAHBLTl0OI,
output
wire
CAHBLTO1OI,
input
CAHBLTII,
input
[
16
:
0
]
CAHBLTI1OI,
input
[
16
:
0
]
CAHBLTl1OI,
input
[
16
:
0
]
CAHBLTOOII,
output
wire
[
31
:
0
]
CAHBLTIOII,
output
reg
CAHBLTlOII,
output
reg
[
2
:
0
]
CAHBLTOIII,
output
reg
CAHBLTIIII,
output
reg
CAHBLTlIII,
output
wire
[
16
:
0
]
CAHBLTOlII,
output
wire
[
16
:
0
]
CAHBLTIlII,
output
reg
CAHBLTllII,
input
[
31
:
0
]
HRDATA_S0,
input
HREADYOUT_S0,
input
[
31
:
0
]
HRDATA_S1,
input
HREADYOUT_S1,
input
[
31
:
0
]
HRDATA_S2,
input
HREADYOUT_S2,
input
[
31
:
0
]
HRDATA_S3,
input
HREADYOUT_S3,
input
[
31
:
0
]
HRDATA_S4,
input
HREADYOUT_S4,
input
[
31
:
0
]
HRDATA_S5,
input
HREADYOUT_S5,
input
[
31
:
0
]
HRDATA_S6,
input
HREADYOUT_S6,
input
[
31
:
0
]
HRDATA_S7,
input
HREADYOUT_S7,
input
[
31
:
0
]
HRDATA_S8,
input
HREADYOUT_S8,
input
[
31
:
0
]
HRDATA_S9,
input
HREADYOUT_S9,
input
[
31
:
0
]
HRDATA_S10,
input
HREADYOUT_S10,
input
[
31
:
0
]
HRDATA_S11,
input
HREADYOUT_S11,
input
[
31
:
0
]
HRDATA_S12,
input
HREADYOUT_S12,
input
[
31
:
0
]
HRDATA_S13,
input
HREADYOUT_S13,
input
[
31
:
0
]
HRDATA_S14,
input
HREADYOUT_S14,
input
[
31
:
0
]
HRDATA_S15,
input
HREADYOUT_S15,
input
[
31
:
0
]
HRDATA_S16,
input
HREADYOUT_S16
)
;
localparam
CAHBLTl0l
=
1
'b
0
;
localparam
CAHBLTO0II
=
1
'b
1
;
localparam
CAHBLTI0II
=
17
'b
0_0000_0000_0000_0000
;
reg
[
31
:
0
]
CAHBLTl0II
;
reg
CAHBLTO1II
;
reg
CAHBLTI1II
;
reg
CAHBLTl1II
;
reg
[
31
:
0
]
CAHBLTOOlI
;
reg
CAHBLTIOlI
;
reg
[
2
:
0
]
CAHBLTlOlI
;
reg
CAHBLTOIlI
;
reg
CAHBLTIIlI
;
reg
CAHBLTlIlI
;
reg
CAHBLTOllI
;
wire
[
16
:
0
]
CAHBLTIllI
;
reg
[
16
:
0
]
CAHBLTlllI
;
reg
[
16
:
0
]
CAHBLTO0lI
;
wire
CAHBLTO0l
;
wire
CAHBLTI0l
;
wire
CAHBLTlll
;
wire
CAHBLTI0lI
;
wire
CAHBLTl0lI
;
wire
CAHBLTO1lI
;
wire
CAHBLTI1lI
;
wire
CAHBLTl1lI
;
wire
CAHBLTOO0I
;
wire
CAHBLTIO0I
;
wire
CAHBLTlO0I
;
wire
CAHBLTOI0I
;
wire
CAHBLTII0I
;
wire
CAHBLTlI0I
;
wire
CAHBLTOl0I
;
wire
CAHBLTIl0I
;
wire
CAHBLTll0I
;
wire
CAHBLTO00I
;
wire
CAHBLTI00I
;
wire
CAHBLTl00I
;
wire
CAHBLTO10I
;
reg
CAHBLTI10I
;
reg
CAHBLTl10I
;
reg
CAHBLTOO1I
;
wire
CAHBLTOO0
;
wire
CAHBLTIO0
;
assign
CAHBLTOO0
=
(
SYNC_RESET
==
1
)
?
1
'b
1
:
HRESETN
;
assign
CAHBLTIO0
=
(
SYNC_RESET
==
1
)
?
HRESETN
:
1
'b
1
;
assign
CAHBLTOlII
=
CAHBLTlllI
[
16
:
0
]
;
assign
CAHBLTIlII
=
CAHBLTO0lI
[
16
:
0
]
;
assign
CAHBLTI0lI
=
(
CAHBLTO0lI
[
0
]
&
(
!
CAHBLTl
[
0
]
)
)
;
assign
CAHBLTl0lI
=
(
CAHBLTO0lI
[
1
]
&
(
!
CAHBLTl
[
1
]
)
)
;
assign
CAHBLTO1lI
=
(
CAHBLTO0lI
[
2
]
&
(
!
CAHBLTl
[
2
]
)
)
;
assign
CAHBLTI1lI
=
(
CAHBLTO0lI
[
3
]
&
(
!
CAHBLTl
[
3
]
)
)
;
assign
CAHBLTl1lI
=
(
CAHBLTO0lI
[
4
]
&
(
!
CAHBLTl
[
4
]
)
)
;
assign
CAHBLTOO0I
=
(
CAHBLTO0lI
[
5
]
&
(
!
CAHBLTl
[
5
]
)
)
;
assign
CAHBLTIO0I
=
(
CAHBLTO0lI
[
6
]
&
(
!
CAHBLTl
[
6
]
)
)
;
assign
CAHBLTlO0I
=
(
CAHBLTO0lI
[
7
]
&
(
!
CAHBLTl
[
7
]
)
)
;
assign
CAHBLTOI0I
=
(
CAHBLTO0lI
[
8
]
&
(
!
CAHBLTl
[
8
]
)
)
;
assign
CAHBLTII0I
=
(
CAHBLTO0lI
[
9
]
&
(
!
CAHBLTl
[
9
]
)
)
;
assign
CAHBLTlI0I
=
(
CAHBLTO0lI
[
10
]
&
(
!
CAHBLTl
[
10
]
)
)
;
assign
CAHBLTOl0I
=
(
CAHBLTO0lI
[
11
]
&
(
!
CAHBLTl
[
11
]
)
)
;
assign
CAHBLTIl0I
=
(
CAHBLTO0lI
[
12
]
&
(
!
CAHBLTl
[
12
]
)
)
;
assign
CAHBLTll0I
=
(
CAHBLTO0lI
[
13
]
&
(
!
CAHBLTl
[
13
]
)
)
;
assign
CAHBLTO00I
=
(
CAHBLTO0lI
[
14
]
&
(
!
CAHBLTl
[
14
]
)
)
;
assign
CAHBLTI00I
=
(
CAHBLTO0lI
[
15
]
&
(
!
CAHBLTl
[
15
]
)
)
;
assign
CAHBLTl00I
=
(
CAHBLTO0lI
[
16
]
&
(
!
CAHBLTl
[
16
]
)
)
;
assign
CAHBLTlll
=
(
CAHBLTI0lI
|
CAHBLTl0lI
|
CAHBLTO1lI
|
CAHBLTI1lI
|
CAHBLTl1lI
|
CAHBLTOO0I
|
CAHBLTIO0I
|
CAHBLTlO0I
|
CAHBLTOI0I
|
CAHBLTII0I
|
CAHBLTlI0I
|
CAHBLTOl0I
|
CAHBLTIl0I
|
CAHBLTll0I
|
CAHBLTO00I
|
CAHBLTI00I
|
CAHBLTl00I
|
CAHBLTl10I
)
;
always
@
(
posedge
HCLK
or
negedge
CAHBLTOO0
)
begin
if
(
(
!
CAHBLTOO0
)
||
(
!
CAHBLTIO0
)
)
begin
CAHBLTOOlI
<=
32
'h
0
;
CAHBLTIOlI
<=
1
'b
0
;
CAHBLTlOlI
<=
3
'b
0
;
CAHBLTOIlI
<=
1
'b
0
;
CAHBLTIIlI
<=
1
'b
0
;
end
else
begin
if
(
CAHBLTl1II
)
begin
CAHBLTOOlI
<=
CAHBLTlIOI
;
CAHBLTIOlI
<=
CAHBLTOlOI
;
CAHBLTlOlI
<=
CAHBLTIlOI
;
CAHBLTOIlI
<=
CAHBLTllOI
;
CAHBLTIIlI
<=
CAHBLTO0OI
;
end
end
end
always
@
(
*
)
begin
if
(
CAHBLTO1II
==
1
'b
0
)
begin
CAHBLTl0II
=
CAHBLTlIOI
;
CAHBLTlOII
=
CAHBLTOlOI
;
CAHBLTOIII
=
CAHBLTIlOI
;
CAHBLTIIII
=
CAHBLTllOI
;
CAHBLTlIII
=
CAHBLTO0OI
;
end
else
begin
CAHBLTl0II
=
CAHBLTOOlI
;
CAHBLTlOII
=
CAHBLTIOlI
;
CAHBLTOIII
=
CAHBLTlOlI
;
CAHBLTIIII
=
CAHBLTOIlI
;
CAHBLTlIII
=
CAHBLTIIlI
;
end
end
CAHBLTO
#
(
.MEMSPACE
(
MEMSPACE
)
,
.HADDR_SHG_CFG
(
HADDR_SHG_CFG
)
,
.CAHBLTI
(
CAHBLTI
)
,
.CAHBLTl
(
CAHBLTl
)
)
CAHBLTIO1I
(
.CAHBLTOI
(
CAHBLTl0II
)
,
.CAHBLTII
(
CAHBLTII
)
,
.CAHBLTlI
(
CAHBLTIllI
[
16
:
0
]
)
,
.CAHBLTOl
(
CAHBLTIOII
[
31
:
0
]
)
,
.CAHBLTIl
(
CAHBLTO10I
)
)
;
always
@
(
*
)
begin
if
(
CAHBLTIIII
)
begin
CAHBLTlllI
=
CAHBLTIllI
;
CAHBLTI10I
=
CAHBLTO10I
;
end
else
begin
CAHBLTlllI
=
CAHBLTI0II
;
CAHBLTI10I
=
1
'b
0
;
end
end
always
@
(
posedge
HCLK
or
negedge
CAHBLTOO0
)
begin
if
(
(
!
CAHBLTOO0
)
||
(
!
CAHBLTIO0
)
)
CAHBLTO0lI
<=
CAHBLTI0II
;
else
if
(
CAHBLTllII
)
CAHBLTO0lI
<=
CAHBLTlllI
;
end
always
@
(
posedge
HCLK
or
negedge
CAHBLTOO0
)
begin
if
(
(
!
CAHBLTOO0
)
||
(
!
CAHBLTIO0
)
)
begin
CAHBLTl10I
<=
1
'b
0
;
end
else
if
(
CAHBLTllII
)
begin
CAHBLTl10I
<=
CAHBLTI10I
;
end
end
always
@
(
*
)
begin
if
(
CAHBLTl10I
)
begin
CAHBLTOO1I
=
CAHBLTO0l
;
CAHBLTI0OI
=
CAHBLTI0l
;
CAHBLTl0OI
=
32
'h
0
;
CAHBLTllII
=
CAHBLTO0l
;
end
else
casez
(
CAHBLTO0lI
[
16
:
0
]
)
17
'b
????????????????1
:
begin
if
(
CAHBLTl
[
0
]
)
begin
CAHBLTOO1I
=
CAHBLTl1OI
[
0
]
;
CAHBLTI0OI
=
CAHBLTOOII
[
0
]
;
CAHBLTl0OI
=
HRDATA_S0
;
CAHBLTllII
=
HREADYOUT_S0
;
end
else
begin
CAHBLTOO1I
=
CAHBLTO0l
;
CAHBLTI0OI
=
CAHBLTI0l
;
CAHBLTl0OI
=
32
'h
0
;
CAHBLTllII
=
CAHBLTO0l
;
end
end
17
'b
???????????????1?
:
begin
if
(
CAHBLTl
[
1
]
)
begin
CAHBLTOO1I
=
CAHBLTl1OI
[
1
]
;
CAHBLTI0OI
=
CAHBLTOOII
[
1
]
;
CAHBLTl0OI
=
HRDATA_S1
;
CAHBLTllII
=
HREADYOUT_S1
;
end
else
begin
CAHBLTOO1I
=
CAHBLTO0l
;
CAHBLTI0OI
=
CAHBLTI0l
;
CAHBLTl0OI
=
32
'h
0
;
CAHBLTllII
=
CAHBLTO0l
;
end
end
17
'b
??????????????1??
:
begin
if
(
CAHBLTl
[
2
]
)
begin
CAHBLTOO1I
=
CAHBLTl1OI
[
2
]
;
CAHBLTI0OI
=
CAHBLTOOII
[
2
]
;
CAHBLTl0OI
=
HRDATA_S2
;
CAHBLTllII
=
HREADYOUT_S2
;
end
else
begin
CAHBLTOO1I
=
CAHBLTO0l
;
CAHBLTI0OI
=
CAHBLTI0l
;
CAHBLTl0OI
=
32
'h
0
;
CAHBLTllII
=
CAHBLTO0l
;
end
end
17
'b
?????????????1???
:
begin
if
(
CAHBLTl
[
3
]
)
begin
CAHBLTOO1I
=
CAHBLTl1OI
[
3
]
;
CAHBLTI0OI
=
CAHBLTOOII
[
3
]
;
CAHBLTl0OI
=
HRDATA_S3
;
CAHBLTllII
=
HREADYOUT_S3
;
end
else
begin
CAHBLTOO1I
=
CAHBLTO0l
;
CAHBLTI0OI
=
CAHBLTI0l
;
CAHBLTl0OI
=
32
'h
0
;
CAHBLTllII
=
CAHBLTO0l
;
end
end
17
'b
????????????1????
:
begin
if
(
CAHBLTl
[
4
]
)
begin
CAHBLTOO1I
=
CAHBLTl1OI
[
4
]
;
CAHBLTI0OI
=
CAHBLTOOII
[
4
]
;
CAHBLTl0OI
=
HRDATA_S4
;
CAHBLTllII
=
HREADYOUT_S4
;
end
else
begin
CAHBLTOO1I
=
CAHBLTO0l
;
CAHBLTI0OI
=
CAHBLTI0l
;
CAHBLTl0OI
=
32
'h
0
;
CAHBLTllII
=
CAHBLTO0l
;
end
end
17
'b
???????????1?????
:
begin
if
(
CAHBLTl
[
5
]
)
begin
CAHBLTOO1I
=
CAHBLTl1OI
[
5
]
;
CAHBLTI0OI
=
CAHBLTOOII
[
5
]
;
CAHBLTl0OI
=
HRDATA_S5
;
CAHBLTllII
=
HREADYOUT_S5
;
end
else
begin
CAHBLTOO1I
=
CAHBLTO0l
;
CAHBLTI0OI
=
CAHBLTI0l
;
CAHBLTl0OI
=
32
'h
0
;
CAHBLTllII
=
CAHBLTO0l
;
end
end
17
'b
??????????1??????
:
begin
if
(
CAHBLTl
[
6
]
)
begin
CAHBLTOO1I
=
CAHBLTl1OI
[
6
]
;
CAHBLTI0OI
=
CAHBLTOOII
[
6
]
;
CAHBLTl0OI
=
HRDATA_S6
;
CAHBLTllII
=
HREADYOUT_S6
;
end
else
begin
CAHBLTOO1I
=
CAHBLTO0l
;
CAHBLTI0OI
=
CAHBLTI0l
;
CAHBLTl0OI
=
32
'h
0
;
CAHBLTllII
=
CAHBLTO0l
;
end
end
17
'b
?????????1???????
:
begin
if
(
CAHBLTl
[
7
]
)
begin
CAHBLTOO1I
=
CAHBLTl1OI
[
7
]
;
CAHBLTI0OI
=
CAHBLTOOII
[
7
]
;
CAHBLTl0OI
=
HRDATA_S7
;
CAHBLTllII
=
HREADYOUT_S7
;
end
else
begin
CAHBLTOO1I
=
CAHBLTO0l
;
CAHBLTI0OI
=
CAHBLTI0l
;
CAHBLTl0OI
=
32
'h
0
;
CAHBLTllII
=
CAHBLTO0l
;
end
end
17
'b
????????1????????
:
begin
if
(
CAHBLTl
[
8
]
)
begin
CAHBLTOO1I
=
CAHBLTl1OI
[
8
]
;
CAHBLTI0OI
=
CAHBLTOOII
[
8
]
;
CAHBLTl0OI
=
HRDATA_S8
;
CAHBLTllII
=
HREADYOUT_S8
;
end
else
begin
CAHBLTOO1I
=
CAHBLTO0l
;
CAHBLTI0OI
=
CAHBLTI0l
;
CAHBLTl0OI
=
32
'h
0
;
CAHBLTllII
=
CAHBLTO0l
;
end
end
17
'b
???????1?????????
:
begin
if
(
CAHBLTl
[
9
]
)
begin
CAHBLTOO1I
=
CAHBLTl1OI
[
9
]
;
CAHBLTI0OI
=
CAHBLTOOII
[
9
]
;
CAHBLTl0OI
=
HRDATA_S9
;
CAHBLTllII
=
HREADYOUT_S9
;
end
else
begin
CAHBLTOO1I
=
CAHBLTO0l
;
CAHBLTI0OI
=
CAHBLTI0l
;
CAHBLTl0OI
=
32
'h
0
;
CAHBLTllII
=
CAHBLTO0l
;
end
end
17
'b
??????1??????????
:
begin
if
(
CAHBLTl
[
10
]
)
begin
CAHBLTOO1I
=
CAHBLTl1OI
[
10
]
;
CAHBLTI0OI
=
CAHBLTOOII
[
10
]
;
CAHBLTl0OI
=
HRDATA_S10
;
CAHBLTllII
=
HREADYOUT_S10
;
end
else
begin
CAHBLTOO1I
=
CAHBLTO0l
;
CAHBLTI0OI
=
CAHBLTI0l
;
CAHBLTl0OI
=
32
'h
0
;
CAHBLTllII
=
CAHBLTO0l
;
end
end
17
'b
?????1???????????
:
begin
if
(
CAHBLTl
[
11
]
)
begin
CAHBLTOO1I
=
CAHBLTl1OI
[
11
]
;
CAHBLTI0OI
=
CAHBLTOOII
[
11
]
;
CAHBLTl0OI
=
HRDATA_S11
;
CAHBLTllII
=
HREADYOUT_S11
;
end
else
begin
CAHBLTOO1I
=
CAHBLTO0l
;
CAHBLTI0OI
=
CAHBLTI0l
;
CAHBLTl0OI
=
32
'h
0
;
CAHBLTllII
=
CAHBLTO0l
;
end
end
17
'b
????1????????????
:
begin
if
(
CAHBLTl
[
12
]
)
begin
CAHBLTOO1I
=
CAHBLTl1OI
[
12
]
;
CAHBLTI0OI
=
CAHBLTOOII
[
12
]
;
CAHBLTl0OI
=
HRDATA_S12
;
CAHBLTllII
=
HREADYOUT_S12
;
end
else
begin
CAHBLTOO1I
=
CAHBLTO0l
;
CAHBLTI0OI
=
CAHBLTI0l
;
CAHBLTl0OI
=
32
'h
0
;
CAHBLTllII
=
CAHBLTO0l
;
end
end
17
'b
???1?????????????
:
begin
if
(
CAHBLTl
[
13
]
)
begin
CAHBLTOO1I
=
CAHBLTl1OI
[
13
]
;
CAHBLTI0OI
=
CAHBLTOOII
[
13
]
;
CAHBLTl0OI
=
HRDATA_S13
;
CAHBLTllII
=
HREADYOUT_S13
;
end
else
begin
CAHBLTOO1I
=
CAHBLTO0l
;
CAHBLTI0OI
=
CAHBLTI0l
;
CAHBLTl0OI
=
32
'h
0
;
CAHBLTllII
=
CAHBLTO0l
;
end
end
17
'b
??1??????????????
:
begin
if
(
CAHBLTl
[
14
]
)
begin
CAHBLTOO1I
=
CAHBLTl1OI
[
14
]
;
CAHBLTI0OI
=
CAHBLTOOII
[
14
]
;
CAHBLTl0OI
=
HRDATA_S14
;
CAHBLTllII
=
HREADYOUT_S14
;
end
else
begin
CAHBLTOO1I
=
CAHBLTO0l
;
CAHBLTI0OI
=
CAHBLTI0l
;
CAHBLTl0OI
=
32
'h
0
;
CAHBLTllII
=
CAHBLTO0l
;
end
end
17
'b
?1???????????????
:
begin
if
(
CAHBLTl
[
15
]
)
begin
CAHBLTOO1I
=
CAHBLTl1OI
[
15
]
;
CAHBLTI0OI
=
CAHBLTOOII
[
15
]
;
CAHBLTl0OI
=
HRDATA_S15
;
CAHBLTllII
=
HREADYOUT_S15
;
end
else
begin
CAHBLTOO1I
=
CAHBLTO0l
;
CAHBLTI0OI
=
CAHBLTI0l
;
CAHBLTl0OI
=
32
'h
0
;
CAHBLTllII
=
CAHBLTO0l
;
end
end
17
'b
1????????????????
:
begin
if
(
CAHBLTl
[
16
]
)
begin
CAHBLTOO1I
=
CAHBLTl1OI
[
16
]
;
CAHBLTI0OI
=
CAHBLTOOII
[
16
]
;
CAHBLTl0OI
=
HRDATA_S16
;
CAHBLTllII
=
HREADYOUT_S16
;
end
else
begin
CAHBLTOO1I
=
CAHBLTO0l
;
CAHBLTI0OI
=
CAHBLTI0l
;
CAHBLTl0OI
=
32
'h
0
;
CAHBLTllII
=
CAHBLTO0l
;
end
end
default
:
begin
CAHBLTOO1I
=
1
'b
1
;
CAHBLTI0OI
=
1
'b
0
;
CAHBLTl0OI
=
32
'h
0
;
CAHBLTllII
=
1
'b
1
;
end
endcase
end
always
@
(
*
)
begin
CAHBLTl1II
=
1
'b
0
;
CAHBLTI1II
=
1
'b
0
;
case
(
CAHBLTlIlI
)
CAHBLTl0l
:
begin
if
(
CAHBLTllOI
&&
CAHBLTO1OI
&&
(
(
CAHBLTIllI
[
0
]
&&
!
CAHBLTI1OI
[
0
]
)
||
(
CAHBLTIllI
[
1
]
&&
!
CAHBLTI1OI
[
1
]
)
||
(
CAHBLTIllI
[
2
]
&&
!
CAHBLTI1OI
[
2
]
)
||
(
CAHBLTIllI
[
3
]
&&
!
CAHBLTI1OI
[
3
]
)
||
(
CAHBLTIllI
[
4
]
&&
!
CAHBLTI1OI
[
4
]
)
||
(
CAHBLTIllI
[
5
]
&&
!
CAHBLTI1OI
[
5
]
)
||
(
CAHBLTIllI
[
6
]
&&
!
CAHBLTI1OI
[
6
]
)
||
(
CAHBLTIllI
[
7
]
&&
!
CAHBLTI1OI
[
7
]
)
||
(
CAHBLTIllI
[
8
]
&&
!
CAHBLTI1OI
[
8
]
)
||
(
CAHBLTIllI
[
9
]
&&
!
CAHBLTI1OI
[
9
]
)
||
(
CAHBLTIllI
[
10
]
&&
!
CAHBLTI1OI
[
10
]
)
||
(
CAHBLTIllI
[
11
]
&&
!
CAHBLTI1OI
[
11
]
)
||
(
CAHBLTIllI
[
12
]
&&
!
CAHBLTI1OI
[
12
]
)
||
(
CAHBLTIllI
[
13
]
&&
!
CAHBLTI1OI
[
13
]
)
||
(
CAHBLTIllI
[
14
]
&&
!
CAHBLTI1OI
[
14
]
)
||
(
CAHBLTIllI
[
15
]
&&
!
CAHBLTI1OI
[
15
]
)
||
(
CAHBLTIllI
[
16
]
&&
!
CAHBLTI1OI
[
16
]
)
)
)
begin
CAHBLTl1II
=
1
'b
1
;
CAHBLTI1II
=
1
'b
1
;
CAHBLTOllI
=
CAHBLTO0II
;
end
else
CAHBLTOllI
=
CAHBLTl0l
;
end
CAHBLTO0II
:
begin
if
(
(
CAHBLTIllI
[
0
]
&&
CAHBLTI1OI
[
0
]
)
||
(
CAHBLTIllI
[
1
]
&&
CAHBLTI1OI
[
1
]
)
||
(
CAHBLTIllI
[
2
]
&&
CAHBLTI1OI
[
2
]
)
||
(
CAHBLTIllI
[
3
]
&&
CAHBLTI1OI
[
3
]
)
||
(
CAHBLTIllI
[
4
]
&&
CAHBLTI1OI
[
4
]
)
||
(
CAHBLTIllI
[
5
]
&&
CAHBLTI1OI
[
5
]
)
||
(
CAHBLTIllI
[
6
]
&&
CAHBLTI1OI
[
6
]
)
||
(
CAHBLTIllI
[
7
]
&&
CAHBLTI1OI
[
7
]
)
||
(
CAHBLTIllI
[
8
]
&&
CAHBLTI1OI
[
8
]
)
||
(
CAHBLTIllI
[
9
]
&&
CAHBLTI1OI
[
9
]
)
||
(
CAHBLTIllI
[
10
]
&&
CAHBLTI1OI
[
10
]
)
||
(
CAHBLTIllI
[
11
]
&&
CAHBLTI1OI
[
11
]
)
||
(
CAHBLTIllI
[
12
]
&&
CAHBLTI1OI
[
12
]
)
||
(
CAHBLTIllI
[
13
]
&&
CAHBLTI1OI
[
13
]
)
||
(
CAHBLTIllI
[
14
]
&&
CAHBLTI1OI
[
14
]
)
||
(
CAHBLTIllI
[
15
]
&&
CAHBLTI1OI
[
15
]
)
||
(
CAHBLTIllI
[
16
]
&&
CAHBLTI1OI
[
16
]
)
)
CAHBLTOllI
=
CAHBLTl0l
;
else
begin
CAHBLTI1II
=
1
'b
1
;
CAHBLTOllI
=
CAHBLTO0II
;
end
end
default
:
CAHBLTOllI
=
CAHBLTl0l
;
endcase
end
always
@
(
posedge
HCLK
or
negedge
CAHBLTOO0
)
begin
if
(
(
!
CAHBLTOO0
)
||
(
!
CAHBLTIO0
)
)
begin
CAHBLTlIlI
<=
CAHBLTl0l
;
CAHBLTO1II
<=
1
'b
0
;
end
else
begin
CAHBLTlIlI
<=
CAHBLTOllI
;
CAHBLTO1II
<=
CAHBLTI1II
;
end
end
CAHBLTIll
#
(
.SYNC_RESET
(
SYNC_RESET
)
)
CAHBLTlO1I
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.CAHBLTlll
(
CAHBLTlll
)
,
.CAHBLTO0l
(
CAHBLTO0l
)
,
.CAHBLTI0l
(
CAHBLTI0l
)
)
;
assign
CAHBLTO1OI
=
CAHBLTOO1I
;
endmodule
