// Actel Corporation Proprietary and Confidential
//  Copyright 2008 Actel Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE ACTEL LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
//  Revision Information:
// Jun09    Revision 4.1
// Aug10    Revision 4.2
// SVN Revision Information:
// SVN $Revision: 8508 $
// SVN $Date: 2009-06-15 16:49:49 -0700 (Mon, 15 Jun 2009) $
`timescale 1ns/1ns
module
CoreUARTapb_C0_CoreUARTapb_C0_0_Tx_async
(
CUARTII
,
CUARTll
,
CUARTlI
,
CUARTl0I
,
CUARTO1I
,
CUARTI1I
,
CUARTlO1
,
CUARTOI1
,
CUARTII1
,
CUARTlI1
,
CUARTOl1
,
CUARTIl1
,
CUARTll1
,
CUARTlll
)
;
parameter
SYNC_RESET
=
0
;
parameter
TX_FIFO
=
0
;
input
CUARTII
;
input
CUARTll
;
input
CUARTlI
;
input
CUARTl0I
;
input
[
7
:
0
]
CUARTO1I
;
input
[
7
:
0
]
CUARTI1I
;
input
CUARTlO1
;
input
CUARTOI1
;
input
CUARTII1
;
input
CUARTlI1
;
input
CUARTOl1
;
output
CUARTIl1
;
wire
CUARTIl1
;
output
CUARTll1
;
output
CUARTlll
;
reg
CUARTll1
;
parameter
CUARTI1ll
=
0
;
parameter
CUARTl1ll
=
1
;
parameter
CUARTOO0l
=
2
;
parameter
CUARTIO0l
=
3
;
parameter
CUARTlO0l
=
4
;
parameter
CUARTOI0l
=
5
;
parameter
CUARTII0l
=
6
;
integer
CUARTlI0l
;
reg
CUARTOl0l
;
reg
[
7
:
0
]
CUARTIl0l
;
reg
[
3
:
0
]
CUARTll0l
;
reg
CUARTO00l
;
wire
CUARTlll
;
reg
CUARTI00l
;
wire
CUARTI1
;
wire
CUARTl1
;
assign
CUARTI1
=
(
SYNC_RESET
==
1
)
?
1
'b
1
:
CUARTlI
;
assign
CUARTl1
=
(
SYNC_RESET
==
1
)
?
CUARTlI
:
1
'b
1
;
always
@
(
posedge
CUARTII
or
negedge
CUARTI1
)
begin
:
CUARTl00l
if
(
(
!
CUARTI1
)
||
(
!
CUARTl1
)
)
begin
CUARTOl0l
<=
1
'b
1
;
end
else
begin
if
(
TX_FIFO
==
1
'b
0
)
begin
if
(
CUARTll
)
begin
if
(
CUARTlI0l
==
CUARTOO0l
)
begin
CUARTOl0l
<=
1
'b
1
;
end
end
if
(
CUARTl0I
)
begin
CUARTOl0l
<=
1
'b
0
;
end
end
else
begin
CUARTOl0l
<=
!
CUARTOI1
;
end
end
end
always
@
(
posedge
CUARTII
or
negedge
CUARTI1
)
begin
:
CUARTO10l
if
(
(
!
CUARTI1
)
||
(
!
CUARTl1
)
)
begin
CUARTlI0l
<=
CUARTI1ll
;
CUARTIl0l
<=
8
'b
0
;
CUARTI00l
<=
1
'b
1
;
end
else
begin
if
(
CUARTll
||
(
CUARTlI0l
==
CUARTI1ll
)
||
(
CUARTlI0l
==
CUARTII0l
)
||
(
CUARTlI0l
==
CUARTl1ll
)
)
begin
CUARTI00l
<=
1
'b
1
;
case
(
CUARTlI0l
)
CUARTI1ll
:
begin
if
(
TX_FIFO
==
1
'b
0
)
begin
if
(
!
CUARTOl0l
)
begin
CUARTlI0l
<=
CUARTl1ll
;
end
else
begin
CUARTlI0l
<=
CUARTI1ll
;
end
end
else
begin
if
(
CUARTlO1
==
1
'b
0
)
begin
CUARTI00l
<=
1
'b
0
;
CUARTlI0l
<=
CUARTII0l
;
end
else
begin
CUARTlI0l
<=
CUARTI1ll
;
CUARTI00l
<=
1
'b
1
;
end
end
end
CUARTl1ll
:
begin
CUARTlI0l
<=
CUARTOO0l
;
end
CUARTOO0l
:
begin
CUARTlI0l
<=
CUARTIO0l
;
if
(
TX_FIFO
==
1
'b
0
)
begin
CUARTIl0l
<=
CUARTO1I
;
end
else
begin
CUARTIl0l
<=
CUARTI1I
;
end
end
CUARTIO0l
:
begin
if
(
CUARTII1
)
begin
if
(
CUARTll0l
==
4
'b
0111
)
begin
if
(
CUARTlI1
)
begin
CUARTlI0l
<=
CUARTlO0l
;
end
else
begin
CUARTlI0l
<=
CUARTOI0l
;
end
end
else
begin
CUARTlI0l
<=
CUARTIO0l
;
end
end
else
begin
if
(
CUARTll0l
==
4
'b
0110
)
begin
if
(
CUARTlI1
)
begin
CUARTlI0l
<=
CUARTlO0l
;
end
else
begin
CUARTlI0l
<=
CUARTOI0l
;
end
end
else
begin
CUARTlI0l
<=
CUARTIO0l
;
end
end
end
CUARTlO0l
:
begin
CUARTlI0l
<=
CUARTOI0l
;
end
CUARTOI0l
:
begin
CUARTlI0l
<=
CUARTI1ll
;
end
CUARTII0l
:
begin
CUARTlI0l
<=
CUARTl1ll
;
end
default
:
begin
CUARTlI0l
<=
CUARTI1ll
;
end
endcase
end
end
end
assign
CUARTlll
=
CUARTI00l
;
always
@
(
posedge
CUARTII
or
negedge
CUARTI1
)
begin
:
CUARTI10l
if
(
(
!
CUARTI1
)
||
(
!
CUARTl1
)
)
begin
CUARTll0l
<=
4
'b
0000
;
end
else
begin
if
(
CUARTll
)
begin
if
(
CUARTlI0l
!=
CUARTIO0l
)
begin
CUARTll0l
<=
4
'b
0000
;
end
else
begin
CUARTll0l
<=
CUARTll0l
+
1
'b
1
;
end
end
end
end
always
@
(
posedge
CUARTII
or
negedge
CUARTI1
)
begin
:
CUARTl10l
if
(
(
!
CUARTI1
)
||
(
!
CUARTl1
)
)
begin
CUARTll1
<=
1
'b
1
;
end
else
begin
if
(
CUARTll
||
(
CUARTlI0l
==
CUARTI1ll
)
||
(
CUARTlI0l
==
CUARTII0l
)
||
(
CUARTlI0l
==
CUARTl1ll
)
)
begin
case
(
CUARTlI0l
)
CUARTI1ll
:
begin
CUARTll1
<=
1
'b
1
;
end
CUARTl1ll
:
begin
CUARTll1
<=
1
'b
1
;
end
CUARTOO0l
:
begin
CUARTll1
<=
1
'b
0
;
end
CUARTIO0l
:
begin
CUARTll1
<=
CUARTIl0l
[
CUARTll0l
]
;
end
CUARTlO0l
:
begin
CUARTll1
<=
CUARTOl1
^
CUARTO00l
;
end
CUARTOI0l
:
begin
CUARTll1
<=
1
'b
1
;
end
default
:
begin
CUARTll1
<=
1
'b
1
;
end
endcase
end
end
end
always
@
(
posedge
CUARTII
or
negedge
CUARTI1
)
begin
:
CUARTOO1l
if
(
(
!
CUARTI1
)
||
(
!
CUARTl1
)
)
begin
CUARTO00l
<=
1
'b
0
;
end
else
begin
if
(
CUARTll
&
CUARTlI1
)
begin
if
(
CUARTlI0l
==
CUARTIO0l
)
begin
CUARTO00l
<=
CUARTO00l
^
CUARTIl0l
[
CUARTll0l
]
;
end
else
begin
CUARTO00l
<=
CUARTO00l
;
end
end
if
(
CUARTlI0l
==
CUARTOI0l
)
begin
CUARTO00l
<=
1
'b
0
;
end
end
end
assign
CUARTIl1
=
CUARTOl0l
;
endmodule
