// Actel Corporation Proprietary and Confidential
// Copyright 2010 Actel Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE ACTEL LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
// SVN Revision Information:
// SVN $Revision: 23120 $
// SVN $Date: 2014-07-17 15:26:23 +0100 (Thu, 17 Jul 2014) $
`timescale 1ns/1ps
module
CAHBLTIll
(
input
HCLK,
input
HRESETN,
input
CAHBLTlll,
output
reg
CAHBLTO0l,
output
reg
CAHBLTI0l
)
;
parameter
SYNC_RESET
=
0
;
localparam
CAHBLTl0l
=
1
'b
0
;
localparam
CAHBLTO1l
=
1
'b
1
;
reg
CAHBLTI1l
;
reg
CAHBLTl1l
;
wire
CAHBLTOO0
;
wire
CAHBLTIO0
;
assign
CAHBLTOO0
=
(
SYNC_RESET
==
1
)
?
1
'b
1
:
HRESETN
;
assign
CAHBLTIO0
=
(
SYNC_RESET
==
1
)
?
HRESETN
:
1
'b
1
;
always
@
(
*
)
begin
CAHBLTO0l
=
1
'b
1
;
CAHBLTI0l
=
1
'b
0
;
case
(
CAHBLTl1l
)
CAHBLTl0l
:
begin
if
(
CAHBLTlll
)
begin
CAHBLTO0l
=
1
'b
0
;
CAHBLTI0l
=
1
'b
1
;
CAHBLTI1l
=
CAHBLTO1l
;
end
else
CAHBLTI1l
=
CAHBLTl0l
;
end
CAHBLTO1l
:
begin
CAHBLTI0l
=
1
'b
1
;
CAHBLTI1l
=
CAHBLTl0l
;
end
default
:
CAHBLTI1l
=
CAHBLTl0l
;
endcase
end
always
@
(
posedge
HCLK
or
negedge
CAHBLTOO0
)
begin
if
(
(
!
CAHBLTOO0
)
||
(
!
CAHBLTIO0
)
)
CAHBLTl1l
<=
CAHBLTl0l
;
else
CAHBLTl1l
<=
CAHBLTI1l
;
end
endmodule
