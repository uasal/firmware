/******************************************************************************

    File Name:  reg_if.v
      Version:  4.0
         Date:  Jul 19th, 2009
  Description:  Register Interface
  
  
  SVN Revision Information:
  SVN $Revision: 11632 $
  SVN $Date: 2009-12-16 15:08:37 -0800 (Wed, 16 Dec 2009) $  
  
  

 COPYRIGHT 2009 BY ACTEL 
 THE INFORMATION CONTAINED IN THIS DOCUMENT IS SUBJECT TO LICENSING RESTRICTIONS 
 FROM ACTEL CORP.  IF YOU ARE NOT IN POSSESSION OF WRITTEN AUTHORIZATION FROM 
 ACTEL FOR USE OF THIS FILE, THEN THE FILE SHOULD BE IMMEDIATELY DESTROYED AND 
 NO BACK-UP OF THE FILE SHOULD BE MADE. 
 
FUNCTIONAL DESCRIPTION: 
Refer to the CorePWM Handbook.
******************************************************************************/
`timescale 1ns/1ns
module
reg_if
#
(
parameter
PWM_NUM
=
8
,
parameter
APB_DWIDTH
=
8
,
parameter
FIXED_PRESCALE_EN
=
0
,
parameter
FIXED_PRESCALE
=
8
,
parameter
FIXED_PERIOD_EN
=
0
,
parameter
FIXED_PERIOD
=
8
,
parameter
DAC_MODE
=
0
,
parameter
SHADOW_REG_EN
=
0
,
parameter
FIXED_PWM_POS_EN
=
0
,
parameter
FIXED_PWM_POSEDGE
=
0
,
parameter
FIXED_PWM_NEG_EN
=
0
,
parameter
FIXED_PWM_NEGEDGE
=
0
)
(
input
PCLK,
input
PRESETN,
input
PSEL,
input
PENABLE,
input
PWRITE,
input
[
5
:
0
]
PADDR,
input
[
APB_DWIDTH
-
1
:
0
]
PWDATA,
output
[
APB_DWIDTH
-
1
:
0
]
CPWMO0,
input
[
APB_DWIDTH
-
1
:
0
]
period_cnt,
input
sync_pulse,
input
[
PWM_NUM
-
1
:
0
]
PWM_STRETCH,
output
[
APB_DWIDTH
-
1
:
0
]
period_out_wire,
output
[
APB_DWIDTH
-
1
:
0
]
prescale_out_wire,
output
[
PWM_NUM
:
1
]
pwm_enable_out_wire,
output
[
PWM_NUM
*
APB_DWIDTH
:
1
]
pwm_posedge_out_wire,
output
[
PWM_NUM
*
APB_DWIDTH
:
1
]
pwm_negedge_out_wire
)
;
wire
[
APB_DWIDTH
-
1
:
0
]
CPWMO01
;
wire
[
APB_DWIDTH
-
1
:
0
]
CPWMI01
;
wire
[
16
:
1
]
CPWMl01
;
wire
[
APB_DWIDTH
-
1
:
0
]
CPWMO11
=
0
;
reg
[
APB_DWIDTH
-
1
:
0
]
CPWMI11
;
reg
[
APB_DWIDTH
-
1
:
0
]
CPWMl11
;
reg
[
PWM_NUM
*
APB_DWIDTH
:
1
]
CPWMOOOI
;
reg
[
PWM_NUM
*
APB_DWIDTH
:
1
]
CPWMIOOI
;
reg
[
APB_DWIDTH
-
1
:
0
]
CPWMlOOI
;
reg
[
APB_DWIDTH
-
1
:
0
]
CPWMOIOI
;
reg
[
APB_DWIDTH
-
1
:
0
]
period_reg
;
reg
[
APB_DWIDTH
-
1
:
0
]
prescale_reg
;
reg
[
8
:
1
]
CPWMIIOI
;
reg
[
16
:
9
]
CPWMlIOI
;
reg
[
16
:
1
]
pwm_enable_reg
;
reg
[
PWM_NUM
*
APB_DWIDTH
:
1
]
CPWMOlOI
;
reg
[
PWM_NUM
*
APB_DWIDTH
:
1
]
CPWMIlOI
;
reg
[
PWM_NUM
*
APB_DWIDTH
:
1
]
pwm_posedge_reg
;
reg
[
PWM_NUM
*
APB_DWIDTH
:
1
]
pwm_negedge_reg
;
reg
CPWMllOI
;
always
@
(
negedge
PRESETN
or
posedge
PCLK
)
begin
if
(
!
PRESETN
)
begin
CPWMlOOI
<=
8
;
CPWMOIOI
<=
8
;
CPWMIIOI
<=
0
;
CPWMlIOI
<=
0
;
end
else
begin
if
(
(
PSEL
==
1
'b
1
)
&&
(
PWRITE
==
1
'b
1
)
&&
(
PENABLE
==
1
'b
1
)
)
begin
case
(
PADDR
)
5
'h
00
:
CPWMlOOI
<=
PWDATA
;
5
'h
01
:
CPWMOIOI
<=
PWDATA
;
5
'h
02
:
CPWMIIOI
<=
PWDATA
[
7
:
0
]
;
5
'h
03
:
CPWMlIOI
<=
PWDATA
[
7
:
0
]
;
endcase
end
end
end
genvar
CPWMO0OI
;
generate
for
(
CPWMO0OI
=
1
;
CPWMO0OI
<=
(
PWM_NUM
)
;
CPWMO0OI
=
CPWMO0OI
+
1
)
begin
:
CPWMI0OI
always
@
(
negedge
PRESETN
or
posedge
PCLK
)
begin
if
(
!
PRESETN
)
begin
CPWMOlOI
[
CPWMO0OI
*
APB_DWIDTH
:
(
CPWMO0OI
-
1
)
*
APB_DWIDTH
+
1
]
<=
0
;
CPWMIlOI
[
CPWMO0OI
*
APB_DWIDTH
:
(
CPWMO0OI
-
1
)
*
APB_DWIDTH
+
1
]
<=
0
;
end
else
begin
if
(
(
PSEL
==
1
'b
1
)
&&
(
PWRITE
==
1
'b
1
)
&&
(
PENABLE
==
1
'b
1
)
)
begin
case
(
PADDR
)
(
2
+
CPWMO0OI
*
2
)
:
begin
CPWMOlOI
[
CPWMO0OI
*
APB_DWIDTH
:
(
CPWMO0OI
-
1
)
*
APB_DWIDTH
+
1
]
<=
PWDATA
;
end
(
3
+
CPWMO0OI
*
2
)
:
CPWMIlOI
[
CPWMO0OI
*
APB_DWIDTH
:
(
CPWMO0OI
-
1
)
*
APB_DWIDTH
+
1
]
<=
PWDATA
;
endcase
end
end
end
end
endgenerate
always
@
(
negedge
PRESETN
or
posedge
PCLK
)
begin
if
(
!
PRESETN
)
begin
CPWMllOI
<=
1
'b
0
;
end
else
begin
if
(
(
PSEL
==
1
'b
1
)
&&
(
PWRITE
==
1
'b
1
)
&&
(
PENABLE
==
1
'b
1
)
)
begin
case
(
PADDR
)
57
:
begin
CPWMllOI
<=
PWDATA
[
0
]
;
end
endcase
end
end
end
genvar
CPWMl0OI
;
generate
for
(
CPWMl0OI
=
1
;
CPWMl0OI
<=
(
PWM_NUM
)
;
CPWMl0OI
=
CPWMl0OI
+
1
)
begin
:
CPWMO1OI
always
@
(
negedge
PRESETN
or
posedge
PCLK
)
begin
if
(
!
PRESETN
)
begin
pwm_posedge_reg
[
CPWMl0OI
*
APB_DWIDTH
:
(
CPWMl0OI
-
1
)
*
APB_DWIDTH
+
1
]
<=
0
;
pwm_negedge_reg
[
CPWMl0OI
*
APB_DWIDTH
:
(
CPWMl0OI
-
1
)
*
APB_DWIDTH
+
1
]
<=
0
;
end
else
begin
if
(
(
period_cnt
>=
period_out_wire
)
&&
(
sync_pulse
)
&&
(
CPWMllOI
==
1
'b
1
)
)
begin
pwm_posedge_reg
[
CPWMl0OI
*
APB_DWIDTH
:
(
CPWMl0OI
-
1
)
*
APB_DWIDTH
+
1
]
<=
CPWMOlOI
[
CPWMl0OI
*
APB_DWIDTH
:
(
CPWMl0OI
-
1
)
*
APB_DWIDTH
+
1
]
;
pwm_negedge_reg
[
CPWMl0OI
*
APB_DWIDTH
:
(
CPWMl0OI
-
1
)
*
APB_DWIDTH
+
1
]
<=
CPWMIlOI
[
CPWMl0OI
*
APB_DWIDTH
:
(
CPWMl0OI
-
1
)
*
APB_DWIDTH
+
1
]
;
end
end
end
end
endgenerate
genvar
CPWMI1OI
;
generate
for
(
CPWMI1OI
=
1
;
CPWMI1OI
<=
(
PWM_NUM
)
;
CPWMI1OI
=
CPWMI1OI
+
1
)
begin
:
CPWMl1OI
always
@*
begin
if
(
SHADOW_REG_EN
[
CPWMI1OI
-
1
]
==
1
)
begin
CPWMOOOI
[
CPWMI1OI
*
APB_DWIDTH
:
(
CPWMI1OI
-
1
)
*
APB_DWIDTH
+
1
]
<=
pwm_posedge_reg
[
CPWMI1OI
*
APB_DWIDTH
:
(
CPWMI1OI
-
1
)
*
APB_DWIDTH
+
1
]
;
CPWMIOOI
[
CPWMI1OI
*
APB_DWIDTH
:
(
CPWMI1OI
-
1
)
*
APB_DWIDTH
+
1
]
<=
pwm_negedge_reg
[
CPWMI1OI
*
APB_DWIDTH
:
(
CPWMI1OI
-
1
)
*
APB_DWIDTH
+
1
]
;
end
else
begin
CPWMOOOI
[
CPWMI1OI
*
APB_DWIDTH
:
(
CPWMI1OI
-
1
)
*
APB_DWIDTH
+
1
]
<=
CPWMOlOI
[
CPWMI1OI
*
APB_DWIDTH
:
(
CPWMI1OI
-
1
)
*
APB_DWIDTH
+
1
]
;
CPWMIOOI
[
CPWMI1OI
*
APB_DWIDTH
:
(
CPWMI1OI
-
1
)
*
APB_DWIDTH
+
1
]
<=
CPWMIlOI
[
CPWMI1OI
*
APB_DWIDTH
:
(
CPWMI1OI
-
1
)
*
APB_DWIDTH
+
1
]
;
end
end
end
endgenerate
genvar
CPWMlO1
;
generate
for
(
CPWMlO1
=
1
;
CPWMlO1
<=
(
PWM_NUM
)
;
CPWMlO1
=
CPWMlO1
+
1
)
begin
:
CPWMOOII
if
(
FIXED_PWM_POS_EN
[
CPWMlO1
-
1
]
==
1
)
begin
assign
pwm_posedge_out_wire
[
CPWMlO1
*
APB_DWIDTH
:
(
CPWMlO1
-
1
)
*
APB_DWIDTH
+
1
]
=
FIXED_PWM_POSEDGE
[
CPWMlO1
*
APB_DWIDTH
-
1
:
(
CPWMlO1
-
1
)
*
APB_DWIDTH
]
;
end
else
begin
assign
pwm_posedge_out_wire
[
CPWMlO1
*
APB_DWIDTH
:
(
CPWMlO1
-
1
)
*
APB_DWIDTH
+
1
]
=
CPWMOOOI
[
CPWMlO1
*
APB_DWIDTH
:
(
CPWMlO1
-
1
)
*
APB_DWIDTH
+
1
]
;
end
end
endgenerate
genvar
CPWMIOII
;
generate
for
(
CPWMIOII
=
1
;
CPWMIOII
<=
(
PWM_NUM
)
;
CPWMIOII
=
CPWMIOII
+
1
)
begin
:
CPWMlOII
if
(
FIXED_PWM_NEG_EN
[
CPWMIOII
-
1
]
==
1
)
begin
assign
pwm_negedge_out_wire
[
CPWMIOII
*
APB_DWIDTH
:
(
CPWMIOII
-
1
)
*
APB_DWIDTH
+
1
]
=
FIXED_PWM_NEGEDGE
[
CPWMIOII
*
APB_DWIDTH
-
1
:
(
CPWMIOII
-
1
)
*
APB_DWIDTH
]
;
end
else
begin
assign
pwm_negedge_out_wire
[
CPWMIOII
*
APB_DWIDTH
:
(
CPWMIOII
-
1
)
*
APB_DWIDTH
+
1
]
=
CPWMIOOI
[
CPWMIOII
*
APB_DWIDTH
:
(
CPWMIOII
-
1
)
*
APB_DWIDTH
+
1
]
;
end
end
endgenerate
always
@
(
negedge
PRESETN
or
posedge
PCLK
)
begin
if
(
!
PRESETN
)
begin
prescale_reg
<=
8
;
period_reg
<=
8
;
pwm_enable_reg
<=
0
;
end
else
begin
if
(
(
period_cnt
>=
period_out_wire
)
&&
(
sync_pulse
)
)
begin
prescale_reg
<=
CPWMlOOI
;
period_reg
<=
CPWMOIOI
;
pwm_enable_reg
<=
{
CPWMlIOI
,
CPWMIIOI
}
;
end
end
end
assign
CPWMl01
=
{
CPWMlIOI
,
CPWMIIOI
}
;
genvar
CPWMOIII
;
generate
for
(
CPWMOIII
=
1
;
CPWMOIII
<=
(
PWM_NUM
)
;
CPWMOIII
=
CPWMOIII
+
1
)
begin
:
CPWMIIII
if
(
SHADOW_REG_EN
[
CPWMOIII
-
1
]
==
1
)
begin
assign
pwm_enable_out_wire
[
CPWMOIII
]
=
pwm_enable_reg
[
CPWMOIII
]
;
end
else
begin
assign
pwm_enable_out_wire
[
CPWMOIII
]
=
CPWMl01
[
CPWMOIII
]
;
end
end
endgenerate
assign
CPWMO01
=
prescale_reg
;
assign
CPWMI01
=
period_reg
;
assign
prescale_out_wire
=
(
FIXED_PRESCALE_EN
==
1
)
?
FIXED_PRESCALE
:
CPWMO01
;
assign
period_out_wire
=
(
FIXED_PERIOD_EN
==
1
)
?
FIXED_PERIOD
:
CPWMI01
;
always
@*
begin
case
(
PADDR
)
0
:
CPWMI11
=
prescale_out_wire
;
1
:
CPWMI11
=
period_out_wire
;
default
:
CPWMI11
=
0
;
endcase
end
generate
if
(
PWM_NUM
==
1
)
begin
:
CPWMIO0
always
@*
begin
case
(
PADDR
)
6
'h
02
:
CPWMl11
=
pwm_enable_out_wire
[
1
]
;
6
'h
03
:
CPWMl11
=
0
;
6
'h
04
:
CPWMl11
=
pwm_posedge_out_wire
[
1
*
APB_DWIDTH
:
0
*
APB_DWIDTH
+
1
]
;
6
'h
05
:
CPWMl11
=
pwm_negedge_out_wire
[
1
*
APB_DWIDTH
:
0
*
APB_DWIDTH
+
1
]
;
6
'h
24
:
CPWMl11
=
PWM_STRETCH
[
PWM_NUM
-
1
:
0
]
;
default
:
CPWMl11
=
0
;
endcase
end
end
endgenerate
generate
if
(
PWM_NUM
==
2
)
begin
:
CPWMlO0
always
@*
begin
case
(
PADDR
)
6
'h
02
:
CPWMl11
=
pwm_enable_out_wire
[
2
:
1
]
;
6
'h
03
:
CPWMl11
=
0
;
6
'h
04
:
CPWMl11
=
pwm_posedge_out_wire
[
1
*
APB_DWIDTH
:
0
*
APB_DWIDTH
+
1
]
;
6
'h
05
:
CPWMl11
=
pwm_negedge_out_wire
[
1
*
APB_DWIDTH
:
0
*
APB_DWIDTH
+
1
]
;
6
'h
06
:
CPWMl11
=
pwm_posedge_out_wire
[
2
*
APB_DWIDTH
:
1
*
APB_DWIDTH
+
1
]
;
6
'h
07
:
CPWMl11
=
pwm_negedge_out_wire
[
2
*
APB_DWIDTH
:
1
*
APB_DWIDTH
+
1
]
;
6
'h
24
:
CPWMl11
=
PWM_STRETCH
[
PWM_NUM
-
1
:
0
]
;
default
:
CPWMl11
=
0
;
endcase
end
end
endgenerate
generate
if
(
PWM_NUM
==
3
)
begin
:
CPWMOI0
always
@*
begin
case
(
PADDR
)
6
'h
02
:
CPWMl11
=
pwm_enable_out_wire
[
3
:
1
]
;
6
'h
03
:
CPWMl11
=
0
;
6
'h
04
:
CPWMl11
=
pwm_posedge_out_wire
[
1
*
APB_DWIDTH
:
0
*
APB_DWIDTH
+
1
]
;
6
'h
05
:
CPWMl11
=
pwm_negedge_out_wire
[
1
*
APB_DWIDTH
:
0
*
APB_DWIDTH
+
1
]
;
6
'h
06
:
CPWMl11
=
pwm_posedge_out_wire
[
2
*
APB_DWIDTH
:
1
*
APB_DWIDTH
+
1
]
;
6
'h
07
:
CPWMl11
=
pwm_negedge_out_wire
[
2
*
APB_DWIDTH
:
1
*
APB_DWIDTH
+
1
]
;
6
'h
08
:
CPWMl11
=
pwm_posedge_out_wire
[
3
*
APB_DWIDTH
:
2
*
APB_DWIDTH
+
1
]
;
6
'h
09
:
CPWMl11
=
pwm_negedge_out_wire
[
3
*
APB_DWIDTH
:
2
*
APB_DWIDTH
+
1
]
;
6
'h
24
:
CPWMl11
=
PWM_STRETCH
[
PWM_NUM
-
1
:
0
]
;
default
:
CPWMl11
=
0
;
endcase
end
end
endgenerate
generate
if
(
PWM_NUM
==
4
)
begin
:
CPWMII0
always
@*
begin
case
(
PADDR
)
6
'h
02
:
CPWMl11
=
pwm_enable_out_wire
[
4
:
1
]
;
6
'h
03
:
CPWMl11
=
0
;
6
'h
04
:
CPWMl11
=
pwm_posedge_out_wire
[
1
*
APB_DWIDTH
:
0
*
APB_DWIDTH
+
1
]
;
6
'h
05
:
CPWMl11
=
pwm_negedge_out_wire
[
1
*
APB_DWIDTH
:
0
*
APB_DWIDTH
+
1
]
;
6
'h
06
:
CPWMl11
=
pwm_posedge_out_wire
[
2
*
APB_DWIDTH
:
1
*
APB_DWIDTH
+
1
]
;
6
'h
07
:
CPWMl11
=
pwm_negedge_out_wire
[
2
*
APB_DWIDTH
:
1
*
APB_DWIDTH
+
1
]
;
6
'h
08
:
CPWMl11
=
pwm_posedge_out_wire
[
3
*
APB_DWIDTH
:
2
*
APB_DWIDTH
+
1
]
;
6
'h
09
:
CPWMl11
=
pwm_negedge_out_wire
[
3
*
APB_DWIDTH
:
2
*
APB_DWIDTH
+
1
]
;
6
'h
0a
:
CPWMl11
=
pwm_posedge_out_wire
[
4
*
APB_DWIDTH
:
3
*
APB_DWIDTH
+
1
]
;
6
'h
0b
:
CPWMl11
=
pwm_negedge_out_wire
[
4
*
APB_DWIDTH
:
3
*
APB_DWIDTH
+
1
]
;
6
'h
24
:
CPWMl11
=
PWM_STRETCH
[
PWM_NUM
-
1
:
0
]
;
default
:
CPWMl11
=
0
;
endcase
end
end
endgenerate
generate
if
(
PWM_NUM
==
5
)
begin
:
CPWMlI0
always
@*
begin
case
(
PADDR
)
6
'h
02
:
CPWMl11
=
pwm_enable_out_wire
[
5
:
1
]
;
6
'h
03
:
CPWMl11
=
0
;
6
'h
04
:
CPWMl11
=
pwm_posedge_out_wire
[
1
*
APB_DWIDTH
:
0
*
APB_DWIDTH
+
1
]
;
6
'h
05
:
CPWMl11
=
pwm_negedge_out_wire
[
1
*
APB_DWIDTH
:
0
*
APB_DWIDTH
+
1
]
;
6
'h
06
:
CPWMl11
=
pwm_posedge_out_wire
[
2
*
APB_DWIDTH
:
1
*
APB_DWIDTH
+
1
]
;
6
'h
07
:
CPWMl11
=
pwm_negedge_out_wire
[
2
*
APB_DWIDTH
:
1
*
APB_DWIDTH
+
1
]
;
6
'h
08
:
CPWMl11
=
pwm_posedge_out_wire
[
3
*
APB_DWIDTH
:
2
*
APB_DWIDTH
+
1
]
;
6
'h
09
:
CPWMl11
=
pwm_negedge_out_wire
[
3
*
APB_DWIDTH
:
2
*
APB_DWIDTH
+
1
]
;
6
'h
0a
:
CPWMl11
=
pwm_posedge_out_wire
[
4
*
APB_DWIDTH
:
3
*
APB_DWIDTH
+
1
]
;
6
'h
0b
:
CPWMl11
=
pwm_negedge_out_wire
[
4
*
APB_DWIDTH
:
3
*
APB_DWIDTH
+
1
]
;
6
'h
0c
:
CPWMl11
=
pwm_posedge_out_wire
[
5
*
APB_DWIDTH
:
4
*
APB_DWIDTH
+
1
]
;
6
'h
0d
:
CPWMl11
=
pwm_negedge_out_wire
[
5
*
APB_DWIDTH
:
4
*
APB_DWIDTH
+
1
]
;
6
'h
24
:
CPWMl11
=
PWM_STRETCH
[
PWM_NUM
-
1
:
0
]
;
default
:
CPWMl11
=
0
;
endcase
end
end
endgenerate
generate
if
(
PWM_NUM
==
6
)
begin
:
CPWMOl0
always
@*
begin
case
(
PADDR
)
6
'h
02
:
CPWMl11
=
pwm_enable_out_wire
[
6
:
1
]
;
6
'h
03
:
CPWMl11
=
0
;
6
'h
04
:
CPWMl11
=
pwm_posedge_out_wire
[
1
*
APB_DWIDTH
:
0
*
APB_DWIDTH
+
1
]
;
6
'h
05
:
CPWMl11
=
pwm_negedge_out_wire
[
1
*
APB_DWIDTH
:
0
*
APB_DWIDTH
+
1
]
;
6
'h
06
:
CPWMl11
=
pwm_posedge_out_wire
[
2
*
APB_DWIDTH
:
1
*
APB_DWIDTH
+
1
]
;
6
'h
07
:
CPWMl11
=
pwm_negedge_out_wire
[
2
*
APB_DWIDTH
:
1
*
APB_DWIDTH
+
1
]
;
6
'h
08
:
CPWMl11
=
pwm_posedge_out_wire
[
3
*
APB_DWIDTH
:
2
*
APB_DWIDTH
+
1
]
;
6
'h
09
:
CPWMl11
=
pwm_negedge_out_wire
[
3
*
APB_DWIDTH
:
2
*
APB_DWIDTH
+
1
]
;
6
'h
0a
:
CPWMl11
=
pwm_posedge_out_wire
[
4
*
APB_DWIDTH
:
3
*
APB_DWIDTH
+
1
]
;
6
'h
0b
:
CPWMl11
=
pwm_negedge_out_wire
[
4
*
APB_DWIDTH
:
3
*
APB_DWIDTH
+
1
]
;
6
'h
0c
:
CPWMl11
=
pwm_posedge_out_wire
[
5
*
APB_DWIDTH
:
4
*
APB_DWIDTH
+
1
]
;
6
'h
0d
:
CPWMl11
=
pwm_negedge_out_wire
[
5
*
APB_DWIDTH
:
4
*
APB_DWIDTH
+
1
]
;
6
'h
0e
:
CPWMl11
=
pwm_posedge_out_wire
[
6
*
APB_DWIDTH
:
5
*
APB_DWIDTH
+
1
]
;
6
'h
0f
:
CPWMl11
=
pwm_negedge_out_wire
[
6
*
APB_DWIDTH
:
5
*
APB_DWIDTH
+
1
]
;
6
'h
24
:
CPWMl11
=
PWM_STRETCH
[
PWM_NUM
-
1
:
0
]
;
default
:
CPWMl11
=
0
;
endcase
end
end
endgenerate
generate
if
(
PWM_NUM
==
7
)
begin
:
CPWMIl0
always
@*
begin
case
(
PADDR
)
6
'h
02
:
CPWMl11
=
pwm_enable_out_wire
[
7
:
1
]
;
6
'h
03
:
CPWMl11
=
0
;
6
'h
04
:
CPWMl11
=
pwm_posedge_out_wire
[
1
*
APB_DWIDTH
:
0
*
APB_DWIDTH
+
1
]
;
6
'h
05
:
CPWMl11
=
pwm_negedge_out_wire
[
1
*
APB_DWIDTH
:
0
*
APB_DWIDTH
+
1
]
;
6
'h
06
:
CPWMl11
=
pwm_posedge_out_wire
[
2
*
APB_DWIDTH
:
1
*
APB_DWIDTH
+
1
]
;
6
'h
07
:
CPWMl11
=
pwm_negedge_out_wire
[
2
*
APB_DWIDTH
:
1
*
APB_DWIDTH
+
1
]
;
6
'h
08
:
CPWMl11
=
pwm_posedge_out_wire
[
3
*
APB_DWIDTH
:
2
*
APB_DWIDTH
+
1
]
;
6
'h
09
:
CPWMl11
=
pwm_negedge_out_wire
[
3
*
APB_DWIDTH
:
2
*
APB_DWIDTH
+
1
]
;
6
'h
0a
:
CPWMl11
=
pwm_posedge_out_wire
[
4
*
APB_DWIDTH
:
3
*
APB_DWIDTH
+
1
]
;
6
'h
0b
:
CPWMl11
=
pwm_negedge_out_wire
[
4
*
APB_DWIDTH
:
3
*
APB_DWIDTH
+
1
]
;
6
'h
0c
:
CPWMl11
=
pwm_posedge_out_wire
[
5
*
APB_DWIDTH
:
4
*
APB_DWIDTH
+
1
]
;
6
'h
0d
:
CPWMl11
=
pwm_negedge_out_wire
[
5
*
APB_DWIDTH
:
4
*
APB_DWIDTH
+
1
]
;
6
'h
0e
:
CPWMl11
=
pwm_posedge_out_wire
[
6
*
APB_DWIDTH
:
5
*
APB_DWIDTH
+
1
]
;
6
'h
0f
:
CPWMl11
=
pwm_negedge_out_wire
[
6
*
APB_DWIDTH
:
5
*
APB_DWIDTH
+
1
]
;
6
'h
10
:
CPWMl11
=
pwm_posedge_out_wire
[
7
*
APB_DWIDTH
:
6
*
APB_DWIDTH
+
1
]
;
6
'h
11
:
CPWMl11
=
pwm_negedge_out_wire
[
7
*
APB_DWIDTH
:
6
*
APB_DWIDTH
+
1
]
;
6
'h
24
:
CPWMl11
=
PWM_STRETCH
[
PWM_NUM
-
1
:
0
]
;
default
:
CPWMl11
=
0
;
endcase
end
end
endgenerate
generate
if
(
PWM_NUM
==
8
)
begin
:
CPWMll0
always
@*
begin
case
(
PADDR
)
6
'h
02
:
CPWMl11
=
pwm_enable_out_wire
[
8
:
1
]
;
6
'h
03
:
CPWMl11
=
0
;
6
'h
04
:
CPWMl11
=
pwm_posedge_out_wire
[
1
*
APB_DWIDTH
:
0
*
APB_DWIDTH
+
1
]
;
6
'h
05
:
CPWMl11
=
pwm_negedge_out_wire
[
1
*
APB_DWIDTH
:
0
*
APB_DWIDTH
+
1
]
;
6
'h
06
:
CPWMl11
=
pwm_posedge_out_wire
[
2
*
APB_DWIDTH
:
1
*
APB_DWIDTH
+
1
]
;
6
'h
07
:
CPWMl11
=
pwm_negedge_out_wire
[
2
*
APB_DWIDTH
:
1
*
APB_DWIDTH
+
1
]
;
6
'h
08
:
CPWMl11
=
pwm_posedge_out_wire
[
3
*
APB_DWIDTH
:
2
*
APB_DWIDTH
+
1
]
;
6
'h
09
:
CPWMl11
=
pwm_negedge_out_wire
[
3
*
APB_DWIDTH
:
2
*
APB_DWIDTH
+
1
]
;
6
'h
0a
:
CPWMl11
=
pwm_posedge_out_wire
[
4
*
APB_DWIDTH
:
3
*
APB_DWIDTH
+
1
]
;
6
'h
0b
:
CPWMl11
=
pwm_negedge_out_wire
[
4
*
APB_DWIDTH
:
3
*
APB_DWIDTH
+
1
]
;
6
'h
0c
:
CPWMl11
=
pwm_posedge_out_wire
[
5
*
APB_DWIDTH
:
4
*
APB_DWIDTH
+
1
]
;
6
'h
0d
:
CPWMl11
=
pwm_negedge_out_wire
[
5
*
APB_DWIDTH
:
4
*
APB_DWIDTH
+
1
]
;
6
'h
0e
:
CPWMl11
=
pwm_posedge_out_wire
[
6
*
APB_DWIDTH
:
5
*
APB_DWIDTH
+
1
]
;
6
'h
0f
:
CPWMl11
=
pwm_negedge_out_wire
[
6
*
APB_DWIDTH
:
5
*
APB_DWIDTH
+
1
]
;
6
'h
10
:
CPWMl11
=
pwm_posedge_out_wire
[
7
*
APB_DWIDTH
:
6
*
APB_DWIDTH
+
1
]
;
6
'h
11
:
CPWMl11
=
pwm_negedge_out_wire
[
7
*
APB_DWIDTH
:
6
*
APB_DWIDTH
+
1
]
;
6
'h
12
:
CPWMl11
=
pwm_posedge_out_wire
[
8
*
APB_DWIDTH
:
7
*
APB_DWIDTH
+
1
]
;
6
'h
13
:
CPWMl11
=
pwm_negedge_out_wire
[
8
*
APB_DWIDTH
:
7
*
APB_DWIDTH
+
1
]
;
6
'h
24
:
CPWMl11
=
PWM_STRETCH
[
PWM_NUM
-
1
:
0
]
;
default
:
CPWMl11
=
0
;
endcase
end
end
endgenerate
generate
if
(
PWM_NUM
==
9
)
begin
:
CPWMO00
always
@*
begin
case
(
PADDR
)
6
'h
02
:
CPWMl11
=
pwm_enable_out_wire
[
8
:
1
]
;
6
'h
03
:
CPWMl11
=
pwm_enable_out_wire
[
9
]
;
6
'h
04
:
CPWMl11
=
pwm_posedge_out_wire
[
1
*
APB_DWIDTH
:
0
*
APB_DWIDTH
+
1
]
;
6
'h
05
:
CPWMl11
=
pwm_negedge_out_wire
[
1
*
APB_DWIDTH
:
0
*
APB_DWIDTH
+
1
]
;
6
'h
06
:
CPWMl11
=
pwm_posedge_out_wire
[
2
*
APB_DWIDTH
:
1
*
APB_DWIDTH
+
1
]
;
6
'h
07
:
CPWMl11
=
pwm_negedge_out_wire
[
2
*
APB_DWIDTH
:
1
*
APB_DWIDTH
+
1
]
;
6
'h
08
:
CPWMl11
=
pwm_posedge_out_wire
[
3
*
APB_DWIDTH
:
2
*
APB_DWIDTH
+
1
]
;
6
'h
09
:
CPWMl11
=
pwm_negedge_out_wire
[
3
*
APB_DWIDTH
:
2
*
APB_DWIDTH
+
1
]
;
6
'h
0a
:
CPWMl11
=
pwm_posedge_out_wire
[
4
*
APB_DWIDTH
:
3
*
APB_DWIDTH
+
1
]
;
6
'h
0b
:
CPWMl11
=
pwm_negedge_out_wire
[
4
*
APB_DWIDTH
:
3
*
APB_DWIDTH
+
1
]
;
6
'h
0c
:
CPWMl11
=
pwm_posedge_out_wire
[
5
*
APB_DWIDTH
:
4
*
APB_DWIDTH
+
1
]
;
6
'h
0d
:
CPWMl11
=
pwm_negedge_out_wire
[
5
*
APB_DWIDTH
:
4
*
APB_DWIDTH
+
1
]
;
6
'h
0e
:
CPWMl11
=
pwm_posedge_out_wire
[
6
*
APB_DWIDTH
:
5
*
APB_DWIDTH
+
1
]
;
6
'h
0f
:
CPWMl11
=
pwm_negedge_out_wire
[
6
*
APB_DWIDTH
:
5
*
APB_DWIDTH
+
1
]
;
6
'h
10
:
CPWMl11
=
pwm_posedge_out_wire
[
7
*
APB_DWIDTH
:
6
*
APB_DWIDTH
+
1
]
;
6
'h
11
:
CPWMl11
=
pwm_negedge_out_wire
[
7
*
APB_DWIDTH
:
6
*
APB_DWIDTH
+
1
]
;
6
'h
12
:
CPWMl11
=
pwm_posedge_out_wire
[
8
*
APB_DWIDTH
:
7
*
APB_DWIDTH
+
1
]
;
6
'h
13
:
CPWMl11
=
pwm_negedge_out_wire
[
8
*
APB_DWIDTH
:
7
*
APB_DWIDTH
+
1
]
;
6
'h
14
:
CPWMl11
=
pwm_posedge_out_wire
[
9
*
APB_DWIDTH
:
8
*
APB_DWIDTH
+
1
]
;
6
'h
15
:
CPWMl11
=
pwm_negedge_out_wire
[
9
*
APB_DWIDTH
:
8
*
APB_DWIDTH
+
1
]
;
6
'h
24
:
CPWMl11
=
PWM_STRETCH
[
PWM_NUM
-
1
:
0
]
;
default
:
CPWMl11
=
0
;
endcase
end
end
endgenerate
generate
if
(
PWM_NUM
==
10
)
begin
:
CPWMI00
always
@*
begin
case
(
PADDR
)
6
'h
02
:
CPWMl11
=
pwm_enable_out_wire
[
8
:
1
]
;
6
'h
03
:
CPWMl11
=
pwm_enable_out_wire
[
10
:
9
]
;
6
'h
04
:
CPWMl11
=
pwm_posedge_out_wire
[
1
*
APB_DWIDTH
:
0
*
APB_DWIDTH
+
1
]
;
6
'h
05
:
CPWMl11
=
pwm_negedge_out_wire
[
1
*
APB_DWIDTH
:
0
*
APB_DWIDTH
+
1
]
;
6
'h
06
:
CPWMl11
=
pwm_posedge_out_wire
[
2
*
APB_DWIDTH
:
1
*
APB_DWIDTH
+
1
]
;
6
'h
07
:
CPWMl11
=
pwm_negedge_out_wire
[
2
*
APB_DWIDTH
:
1
*
APB_DWIDTH
+
1
]
;
6
'h
08
:
CPWMl11
=
pwm_posedge_out_wire
[
3
*
APB_DWIDTH
:
2
*
APB_DWIDTH
+
1
]
;
6
'h
09
:
CPWMl11
=
pwm_negedge_out_wire
[
3
*
APB_DWIDTH
:
2
*
APB_DWIDTH
+
1
]
;
6
'h
0a
:
CPWMl11
=
pwm_posedge_out_wire
[
4
*
APB_DWIDTH
:
3
*
APB_DWIDTH
+
1
]
;
6
'h
0b
:
CPWMl11
=
pwm_negedge_out_wire
[
4
*
APB_DWIDTH
:
3
*
APB_DWIDTH
+
1
]
;
6
'h
0c
:
CPWMl11
=
pwm_posedge_out_wire
[
5
*
APB_DWIDTH
:
4
*
APB_DWIDTH
+
1
]
;
6
'h
0d
:
CPWMl11
=
pwm_negedge_out_wire
[
5
*
APB_DWIDTH
:
4
*
APB_DWIDTH
+
1
]
;
6
'h
0e
:
CPWMl11
=
pwm_posedge_out_wire
[
6
*
APB_DWIDTH
:
5
*
APB_DWIDTH
+
1
]
;
6
'h
0f
:
CPWMl11
=
pwm_negedge_out_wire
[
6
*
APB_DWIDTH
:
5
*
APB_DWIDTH
+
1
]
;
6
'h
10
:
CPWMl11
=
pwm_posedge_out_wire
[
7
*
APB_DWIDTH
:
6
*
APB_DWIDTH
+
1
]
;
6
'h
11
:
CPWMl11
=
pwm_negedge_out_wire
[
7
*
APB_DWIDTH
:
6
*
APB_DWIDTH
+
1
]
;
6
'h
12
:
CPWMl11
=
pwm_posedge_out_wire
[
8
*
APB_DWIDTH
:
7
*
APB_DWIDTH
+
1
]
;
6
'h
13
:
CPWMl11
=
pwm_negedge_out_wire
[
8
*
APB_DWIDTH
:
7
*
APB_DWIDTH
+
1
]
;
6
'h
14
:
CPWMl11
=
pwm_posedge_out_wire
[
9
*
APB_DWIDTH
:
8
*
APB_DWIDTH
+
1
]
;
6
'h
15
:
CPWMl11
=
pwm_negedge_out_wire
[
9
*
APB_DWIDTH
:
8
*
APB_DWIDTH
+
1
]
;
6
'h
16
:
CPWMl11
=
pwm_posedge_out_wire
[
10
*
APB_DWIDTH
:
9
*
APB_DWIDTH
+
1
]
;
6
'h
17
:
CPWMl11
=
pwm_negedge_out_wire
[
10
*
APB_DWIDTH
:
9
*
APB_DWIDTH
+
1
]
;
6
'h
24
:
CPWMl11
=
PWM_STRETCH
[
PWM_NUM
-
1
:
0
]
;
default
:
CPWMl11
=
0
;
endcase
end
end
endgenerate
generate
if
(
PWM_NUM
==
11
)
begin
:
CPWMl00
always
@*
begin
case
(
PADDR
)
6
'h
02
:
CPWMl11
=
pwm_enable_out_wire
[
8
:
1
]
;
6
'h
03
:
CPWMl11
=
pwm_enable_out_wire
[
11
:
9
]
;
6
'h
04
:
CPWMl11
=
pwm_posedge_out_wire
[
1
*
APB_DWIDTH
:
0
*
APB_DWIDTH
+
1
]
;
6
'h
05
:
CPWMl11
=
pwm_negedge_out_wire
[
1
*
APB_DWIDTH
:
0
*
APB_DWIDTH
+
1
]
;
6
'h
06
:
CPWMl11
=
pwm_posedge_out_wire
[
2
*
APB_DWIDTH
:
1
*
APB_DWIDTH
+
1
]
;
6
'h
07
:
CPWMl11
=
pwm_negedge_out_wire
[
2
*
APB_DWIDTH
:
1
*
APB_DWIDTH
+
1
]
;
6
'h
08
:
CPWMl11
=
pwm_posedge_out_wire
[
3
*
APB_DWIDTH
:
2
*
APB_DWIDTH
+
1
]
;
6
'h
09
:
CPWMl11
=
pwm_negedge_out_wire
[
3
*
APB_DWIDTH
:
2
*
APB_DWIDTH
+
1
]
;
6
'h
0a
:
CPWMl11
=
pwm_posedge_out_wire
[
4
*
APB_DWIDTH
:
3
*
APB_DWIDTH
+
1
]
;
6
'h
0b
:
CPWMl11
=
pwm_negedge_out_wire
[
4
*
APB_DWIDTH
:
3
*
APB_DWIDTH
+
1
]
;
6
'h
0c
:
CPWMl11
=
pwm_posedge_out_wire
[
5
*
APB_DWIDTH
:
4
*
APB_DWIDTH
+
1
]
;
6
'h
0d
:
CPWMl11
=
pwm_negedge_out_wire
[
5
*
APB_DWIDTH
:
4
*
APB_DWIDTH
+
1
]
;
6
'h
0e
:
CPWMl11
=
pwm_posedge_out_wire
[
6
*
APB_DWIDTH
:
5
*
APB_DWIDTH
+
1
]
;
6
'h
0f
:
CPWMl11
=
pwm_negedge_out_wire
[
6
*
APB_DWIDTH
:
5
*
APB_DWIDTH
+
1
]
;
6
'h
10
:
CPWMl11
=
pwm_posedge_out_wire
[
7
*
APB_DWIDTH
:
6
*
APB_DWIDTH
+
1
]
;
6
'h
11
:
CPWMl11
=
pwm_negedge_out_wire
[
7
*
APB_DWIDTH
:
6
*
APB_DWIDTH
+
1
]
;
6
'h
12
:
CPWMl11
=
pwm_posedge_out_wire
[
8
*
APB_DWIDTH
:
7
*
APB_DWIDTH
+
1
]
;
6
'h
13
:
CPWMl11
=
pwm_negedge_out_wire
[
8
*
APB_DWIDTH
:
7
*
APB_DWIDTH
+
1
]
;
6
'h
14
:
CPWMl11
=
pwm_posedge_out_wire
[
9
*
APB_DWIDTH
:
8
*
APB_DWIDTH
+
1
]
;
6
'h
15
:
CPWMl11
=
pwm_negedge_out_wire
[
9
*
APB_DWIDTH
:
8
*
APB_DWIDTH
+
1
]
;
6
'h
16
:
CPWMl11
=
pwm_posedge_out_wire
[
10
*
APB_DWIDTH
:
9
*
APB_DWIDTH
+
1
]
;
6
'h
17
:
CPWMl11
=
pwm_negedge_out_wire
[
10
*
APB_DWIDTH
:
9
*
APB_DWIDTH
+
1
]
;
6
'h
18
:
CPWMl11
=
pwm_posedge_out_wire
[
11
*
APB_DWIDTH
:
10
*
APB_DWIDTH
+
1
]
;
6
'h
19
:
CPWMl11
=
pwm_negedge_out_wire
[
11
*
APB_DWIDTH
:
10
*
APB_DWIDTH
+
1
]
;
6
'h
24
:
CPWMl11
=
PWM_STRETCH
[
PWM_NUM
-
1
:
0
]
;
default
:
CPWMl11
=
0
;
endcase
end
end
endgenerate
generate
if
(
PWM_NUM
==
12
)
begin
:
CPWMO10
always
@*
begin
case
(
PADDR
)
6
'h
02
:
CPWMl11
=
pwm_enable_out_wire
[
8
:
1
]
;
6
'h
03
:
CPWMl11
=
pwm_enable_out_wire
[
12
:
9
]
;
6
'h
04
:
CPWMl11
=
pwm_posedge_out_wire
[
1
*
APB_DWIDTH
:
0
*
APB_DWIDTH
+
1
]
;
6
'h
05
:
CPWMl11
=
pwm_negedge_out_wire
[
1
*
APB_DWIDTH
:
0
*
APB_DWIDTH
+
1
]
;
6
'h
06
:
CPWMl11
=
pwm_posedge_out_wire
[
2
*
APB_DWIDTH
:
1
*
APB_DWIDTH
+
1
]
;
6
'h
07
:
CPWMl11
=
pwm_negedge_out_wire
[
2
*
APB_DWIDTH
:
1
*
APB_DWIDTH
+
1
]
;
6
'h
08
:
CPWMl11
=
pwm_posedge_out_wire
[
3
*
APB_DWIDTH
:
2
*
APB_DWIDTH
+
1
]
;
6
'h
09
:
CPWMl11
=
pwm_negedge_out_wire
[
3
*
APB_DWIDTH
:
2
*
APB_DWIDTH
+
1
]
;
6
'h
0a
:
CPWMl11
=
pwm_posedge_out_wire
[
4
*
APB_DWIDTH
:
3
*
APB_DWIDTH
+
1
]
;
6
'h
0b
:
CPWMl11
=
pwm_negedge_out_wire
[
4
*
APB_DWIDTH
:
3
*
APB_DWIDTH
+
1
]
;
6
'h
0c
:
CPWMl11
=
pwm_posedge_out_wire
[
5
*
APB_DWIDTH
:
4
*
APB_DWIDTH
+
1
]
;
6
'h
0d
:
CPWMl11
=
pwm_negedge_out_wire
[
5
*
APB_DWIDTH
:
4
*
APB_DWIDTH
+
1
]
;
6
'h
0e
:
CPWMl11
=
pwm_posedge_out_wire
[
6
*
APB_DWIDTH
:
5
*
APB_DWIDTH
+
1
]
;
6
'h
0f
:
CPWMl11
=
pwm_negedge_out_wire
[
6
*
APB_DWIDTH
:
5
*
APB_DWIDTH
+
1
]
;
6
'h
10
:
CPWMl11
=
pwm_posedge_out_wire
[
7
*
APB_DWIDTH
:
6
*
APB_DWIDTH
+
1
]
;
6
'h
11
:
CPWMl11
=
pwm_negedge_out_wire
[
7
*
APB_DWIDTH
:
6
*
APB_DWIDTH
+
1
]
;
6
'h
12
:
CPWMl11
=
pwm_posedge_out_wire
[
8
*
APB_DWIDTH
:
7
*
APB_DWIDTH
+
1
]
;
6
'h
13
:
CPWMl11
=
pwm_negedge_out_wire
[
8
*
APB_DWIDTH
:
7
*
APB_DWIDTH
+
1
]
;
6
'h
14
:
CPWMl11
=
pwm_posedge_out_wire
[
9
*
APB_DWIDTH
:
8
*
APB_DWIDTH
+
1
]
;
6
'h
15
:
CPWMl11
=
pwm_negedge_out_wire
[
9
*
APB_DWIDTH
:
8
*
APB_DWIDTH
+
1
]
;
6
'h
16
:
CPWMl11
=
pwm_posedge_out_wire
[
10
*
APB_DWIDTH
:
9
*
APB_DWIDTH
+
1
]
;
6
'h
17
:
CPWMl11
=
pwm_negedge_out_wire
[
10
*
APB_DWIDTH
:
9
*
APB_DWIDTH
+
1
]
;
6
'h
18
:
CPWMl11
=
pwm_posedge_out_wire
[
11
*
APB_DWIDTH
:
10
*
APB_DWIDTH
+
1
]
;
6
'h
19
:
CPWMl11
=
pwm_negedge_out_wire
[
11
*
APB_DWIDTH
:
10
*
APB_DWIDTH
+
1
]
;
6
'h
1a
:
CPWMl11
=
pwm_posedge_out_wire
[
12
*
APB_DWIDTH
:
11
*
APB_DWIDTH
+
1
]
;
6
'h
1b
:
CPWMl11
=
pwm_negedge_out_wire
[
12
*
APB_DWIDTH
:
11
*
APB_DWIDTH
+
1
]
;
6
'h
24
:
CPWMl11
=
PWM_STRETCH
[
PWM_NUM
-
1
:
0
]
;
default
:
CPWMl11
=
0
;
endcase
end
end
endgenerate
generate
if
(
PWM_NUM
==
13
)
begin
:
CPWMI10
always
@*
begin
case
(
PADDR
)
6
'h
02
:
CPWMl11
=
pwm_enable_out_wire
[
8
:
1
]
;
6
'h
03
:
CPWMl11
=
pwm_enable_out_wire
[
13
:
9
]
;
6
'h
04
:
CPWMl11
=
pwm_posedge_out_wire
[
1
*
APB_DWIDTH
:
0
*
APB_DWIDTH
+
1
]
;
6
'h
05
:
CPWMl11
=
pwm_negedge_out_wire
[
1
*
APB_DWIDTH
:
0
*
APB_DWIDTH
+
1
]
;
6
'h
06
:
CPWMl11
=
pwm_posedge_out_wire
[
2
*
APB_DWIDTH
:
1
*
APB_DWIDTH
+
1
]
;
6
'h
07
:
CPWMl11
=
pwm_negedge_out_wire
[
2
*
APB_DWIDTH
:
1
*
APB_DWIDTH
+
1
]
;
6
'h
08
:
CPWMl11
=
pwm_posedge_out_wire
[
3
*
APB_DWIDTH
:
2
*
APB_DWIDTH
+
1
]
;
6
'h
09
:
CPWMl11
=
pwm_negedge_out_wire
[
3
*
APB_DWIDTH
:
2
*
APB_DWIDTH
+
1
]
;
6
'h
0a
:
CPWMl11
=
pwm_posedge_out_wire
[
4
*
APB_DWIDTH
:
3
*
APB_DWIDTH
+
1
]
;
6
'h
0b
:
CPWMl11
=
pwm_negedge_out_wire
[
4
*
APB_DWIDTH
:
3
*
APB_DWIDTH
+
1
]
;
6
'h
0c
:
CPWMl11
=
pwm_posedge_out_wire
[
5
*
APB_DWIDTH
:
4
*
APB_DWIDTH
+
1
]
;
6
'h
0d
:
CPWMl11
=
pwm_negedge_out_wire
[
5
*
APB_DWIDTH
:
4
*
APB_DWIDTH
+
1
]
;
6
'h
0e
:
CPWMl11
=
pwm_posedge_out_wire
[
6
*
APB_DWIDTH
:
5
*
APB_DWIDTH
+
1
]
;
6
'h
0f
:
CPWMl11
=
pwm_negedge_out_wire
[
6
*
APB_DWIDTH
:
5
*
APB_DWIDTH
+
1
]
;
6
'h
10
:
CPWMl11
=
pwm_posedge_out_wire
[
7
*
APB_DWIDTH
:
6
*
APB_DWIDTH
+
1
]
;
6
'h
11
:
CPWMl11
=
pwm_negedge_out_wire
[
7
*
APB_DWIDTH
:
6
*
APB_DWIDTH
+
1
]
;
6
'h
12
:
CPWMl11
=
pwm_posedge_out_wire
[
8
*
APB_DWIDTH
:
7
*
APB_DWIDTH
+
1
]
;
6
'h
13
:
CPWMl11
=
pwm_negedge_out_wire
[
8
*
APB_DWIDTH
:
7
*
APB_DWIDTH
+
1
]
;
6
'h
14
:
CPWMl11
=
pwm_posedge_out_wire
[
9
*
APB_DWIDTH
:
8
*
APB_DWIDTH
+
1
]
;
6
'h
15
:
CPWMl11
=
pwm_negedge_out_wire
[
9
*
APB_DWIDTH
:
8
*
APB_DWIDTH
+
1
]
;
6
'h
16
:
CPWMl11
=
pwm_posedge_out_wire
[
10
*
APB_DWIDTH
:
9
*
APB_DWIDTH
+
1
]
;
6
'h
17
:
CPWMl11
=
pwm_negedge_out_wire
[
10
*
APB_DWIDTH
:
9
*
APB_DWIDTH
+
1
]
;
6
'h
18
:
CPWMl11
=
pwm_posedge_out_wire
[
11
*
APB_DWIDTH
:
10
*
APB_DWIDTH
+
1
]
;
6
'h
19
:
CPWMl11
=
pwm_negedge_out_wire
[
11
*
APB_DWIDTH
:
10
*
APB_DWIDTH
+
1
]
;
6
'h
1a
:
CPWMl11
=
pwm_posedge_out_wire
[
12
*
APB_DWIDTH
:
11
*
APB_DWIDTH
+
1
]
;
6
'h
1b
:
CPWMl11
=
pwm_negedge_out_wire
[
12
*
APB_DWIDTH
:
11
*
APB_DWIDTH
+
1
]
;
6
'h
1c
:
CPWMl11
=
pwm_posedge_out_wire
[
13
*
APB_DWIDTH
:
12
*
APB_DWIDTH
+
1
]
;
6
'h
1d
:
CPWMl11
=
pwm_negedge_out_wire
[
13
*
APB_DWIDTH
:
12
*
APB_DWIDTH
+
1
]
;
6
'h
24
:
CPWMl11
=
PWM_STRETCH
[
PWM_NUM
-
1
:
0
]
;
default
:
CPWMl11
=
0
;
endcase
end
end
endgenerate
generate
if
(
PWM_NUM
==
14
)
begin
:
CPWMl10
always
@*
begin
case
(
PADDR
)
6
'h
02
:
CPWMl11
=
pwm_enable_out_wire
[
8
:
1
]
;
6
'h
03
:
CPWMl11
=
pwm_enable_out_wire
[
14
:
9
]
;
6
'h
04
:
CPWMl11
=
pwm_posedge_out_wire
[
1
*
APB_DWIDTH
:
0
*
APB_DWIDTH
+
1
]
;
6
'h
05
:
CPWMl11
=
pwm_negedge_out_wire
[
1
*
APB_DWIDTH
:
0
*
APB_DWIDTH
+
1
]
;
6
'h
06
:
CPWMl11
=
pwm_posedge_out_wire
[
2
*
APB_DWIDTH
:
1
*
APB_DWIDTH
+
1
]
;
6
'h
07
:
CPWMl11
=
pwm_negedge_out_wire
[
2
*
APB_DWIDTH
:
1
*
APB_DWIDTH
+
1
]
;
6
'h
08
:
CPWMl11
=
pwm_posedge_out_wire
[
3
*
APB_DWIDTH
:
2
*
APB_DWIDTH
+
1
]
;
6
'h
09
:
CPWMl11
=
pwm_negedge_out_wire
[
3
*
APB_DWIDTH
:
2
*
APB_DWIDTH
+
1
]
;
6
'h
0a
:
CPWMl11
=
pwm_posedge_out_wire
[
4
*
APB_DWIDTH
:
3
*
APB_DWIDTH
+
1
]
;
6
'h
0b
:
CPWMl11
=
pwm_negedge_out_wire
[
4
*
APB_DWIDTH
:
3
*
APB_DWIDTH
+
1
]
;
6
'h
0c
:
CPWMl11
=
pwm_posedge_out_wire
[
5
*
APB_DWIDTH
:
4
*
APB_DWIDTH
+
1
]
;
6
'h
0d
:
CPWMl11
=
pwm_negedge_out_wire
[
5
*
APB_DWIDTH
:
4
*
APB_DWIDTH
+
1
]
;
6
'h
0e
:
CPWMl11
=
pwm_posedge_out_wire
[
6
*
APB_DWIDTH
:
5
*
APB_DWIDTH
+
1
]
;
6
'h
0f
:
CPWMl11
=
pwm_negedge_out_wire
[
6
*
APB_DWIDTH
:
5
*
APB_DWIDTH
+
1
]
;
6
'h
10
:
CPWMl11
=
pwm_posedge_out_wire
[
7
*
APB_DWIDTH
:
6
*
APB_DWIDTH
+
1
]
;
6
'h
11
:
CPWMl11
=
pwm_negedge_out_wire
[
7
*
APB_DWIDTH
:
6
*
APB_DWIDTH
+
1
]
;
6
'h
12
:
CPWMl11
=
pwm_posedge_out_wire
[
8
*
APB_DWIDTH
:
7
*
APB_DWIDTH
+
1
]
;
6
'h
13
:
CPWMl11
=
pwm_negedge_out_wire
[
8
*
APB_DWIDTH
:
7
*
APB_DWIDTH
+
1
]
;
6
'h
14
:
CPWMl11
=
pwm_posedge_out_wire
[
9
*
APB_DWIDTH
:
8
*
APB_DWIDTH
+
1
]
;
6
'h
15
:
CPWMl11
=
pwm_negedge_out_wire
[
9
*
APB_DWIDTH
:
8
*
APB_DWIDTH
+
1
]
;
6
'h
16
:
CPWMl11
=
pwm_posedge_out_wire
[
10
*
APB_DWIDTH
:
9
*
APB_DWIDTH
+
1
]
;
6
'h
17
:
CPWMl11
=
pwm_negedge_out_wire
[
10
*
APB_DWIDTH
:
9
*
APB_DWIDTH
+
1
]
;
6
'h
18
:
CPWMl11
=
pwm_posedge_out_wire
[
11
*
APB_DWIDTH
:
10
*
APB_DWIDTH
+
1
]
;
6
'h
19
:
CPWMl11
=
pwm_negedge_out_wire
[
11
*
APB_DWIDTH
:
10
*
APB_DWIDTH
+
1
]
;
6
'h
1a
:
CPWMl11
=
pwm_posedge_out_wire
[
12
*
APB_DWIDTH
:
11
*
APB_DWIDTH
+
1
]
;
6
'h
1b
:
CPWMl11
=
pwm_negedge_out_wire
[
12
*
APB_DWIDTH
:
11
*
APB_DWIDTH
+
1
]
;
6
'h
1c
:
CPWMl11
=
pwm_posedge_out_wire
[
13
*
APB_DWIDTH
:
12
*
APB_DWIDTH
+
1
]
;
6
'h
1d
:
CPWMl11
=
pwm_negedge_out_wire
[
13
*
APB_DWIDTH
:
12
*
APB_DWIDTH
+
1
]
;
6
'h
1e
:
CPWMl11
=
pwm_posedge_out_wire
[
14
*
APB_DWIDTH
:
13
*
APB_DWIDTH
+
1
]
;
6
'h
1f
:
CPWMl11
=
pwm_negedge_out_wire
[
14
*
APB_DWIDTH
:
13
*
APB_DWIDTH
+
1
]
;
6
'h
24
:
CPWMl11
=
PWM_STRETCH
[
PWM_NUM
-
1
:
0
]
;
default
:
CPWMl11
=
0
;
endcase
end
end
endgenerate
generate
if
(
PWM_NUM
==
15
)
begin
:
CPWMOO1
always
@*
begin
case
(
PADDR
)
6
'h
02
:
CPWMl11
=
pwm_enable_out_wire
[
8
:
1
]
;
6
'h
03
:
CPWMl11
=
pwm_enable_out_wire
[
15
:
9
]
;
6
'h
04
:
CPWMl11
=
pwm_posedge_out_wire
[
1
*
APB_DWIDTH
:
0
*
APB_DWIDTH
+
1
]
;
6
'h
05
:
CPWMl11
=
pwm_negedge_out_wire
[
1
*
APB_DWIDTH
:
0
*
APB_DWIDTH
+
1
]
;
6
'h
06
:
CPWMl11
=
pwm_posedge_out_wire
[
2
*
APB_DWIDTH
:
1
*
APB_DWIDTH
+
1
]
;
6
'h
07
:
CPWMl11
=
pwm_negedge_out_wire
[
2
*
APB_DWIDTH
:
1
*
APB_DWIDTH
+
1
]
;
6
'h
08
:
CPWMl11
=
pwm_posedge_out_wire
[
3
*
APB_DWIDTH
:
2
*
APB_DWIDTH
+
1
]
;
6
'h
09
:
CPWMl11
=
pwm_negedge_out_wire
[
3
*
APB_DWIDTH
:
2
*
APB_DWIDTH
+
1
]
;
6
'h
0a
:
CPWMl11
=
pwm_posedge_out_wire
[
4
*
APB_DWIDTH
:
3
*
APB_DWIDTH
+
1
]
;
6
'h
0b
:
CPWMl11
=
pwm_negedge_out_wire
[
4
*
APB_DWIDTH
:
3
*
APB_DWIDTH
+
1
]
;
6
'h
0c
:
CPWMl11
=
pwm_posedge_out_wire
[
5
*
APB_DWIDTH
:
4
*
APB_DWIDTH
+
1
]
;
6
'h
0d
:
CPWMl11
=
pwm_negedge_out_wire
[
5
*
APB_DWIDTH
:
4
*
APB_DWIDTH
+
1
]
;
6
'h
0e
:
CPWMl11
=
pwm_posedge_out_wire
[
6
*
APB_DWIDTH
:
5
*
APB_DWIDTH
+
1
]
;
6
'h
0f
:
CPWMl11
=
pwm_negedge_out_wire
[
6
*
APB_DWIDTH
:
5
*
APB_DWIDTH
+
1
]
;
6
'h
10
:
CPWMl11
=
pwm_posedge_out_wire
[
7
*
APB_DWIDTH
:
6
*
APB_DWIDTH
+
1
]
;
6
'h
11
:
CPWMl11
=
pwm_negedge_out_wire
[
7
*
APB_DWIDTH
:
6
*
APB_DWIDTH
+
1
]
;
6
'h
12
:
CPWMl11
=
pwm_posedge_out_wire
[
8
*
APB_DWIDTH
:
7
*
APB_DWIDTH
+
1
]
;
6
'h
13
:
CPWMl11
=
pwm_negedge_out_wire
[
8
*
APB_DWIDTH
:
7
*
APB_DWIDTH
+
1
]
;
6
'h
14
:
CPWMl11
=
pwm_posedge_out_wire
[
9
*
APB_DWIDTH
:
8
*
APB_DWIDTH
+
1
]
;
6
'h
15
:
CPWMl11
=
pwm_negedge_out_wire
[
9
*
APB_DWIDTH
:
8
*
APB_DWIDTH
+
1
]
;
6
'h
16
:
CPWMl11
=
pwm_posedge_out_wire
[
10
*
APB_DWIDTH
:
9
*
APB_DWIDTH
+
1
]
;
6
'h
17
:
CPWMl11
=
pwm_negedge_out_wire
[
10
*
APB_DWIDTH
:
9
*
APB_DWIDTH
+
1
]
;
6
'h
18
:
CPWMl11
=
pwm_posedge_out_wire
[
11
*
APB_DWIDTH
:
10
*
APB_DWIDTH
+
1
]
;
6
'h
19
:
CPWMl11
=
pwm_negedge_out_wire
[
11
*
APB_DWIDTH
:
10
*
APB_DWIDTH
+
1
]
;
6
'h
1a
:
CPWMl11
=
pwm_posedge_out_wire
[
12
*
APB_DWIDTH
:
11
*
APB_DWIDTH
+
1
]
;
6
'h
1b
:
CPWMl11
=
pwm_negedge_out_wire
[
12
*
APB_DWIDTH
:
11
*
APB_DWIDTH
+
1
]
;
6
'h
1c
:
CPWMl11
=
pwm_posedge_out_wire
[
13
*
APB_DWIDTH
:
12
*
APB_DWIDTH
+
1
]
;
6
'h
1d
:
CPWMl11
=
pwm_negedge_out_wire
[
13
*
APB_DWIDTH
:
12
*
APB_DWIDTH
+
1
]
;
6
'h
1e
:
CPWMl11
=
pwm_posedge_out_wire
[
14
*
APB_DWIDTH
:
13
*
APB_DWIDTH
+
1
]
;
6
'h
1f
:
CPWMl11
=
pwm_negedge_out_wire
[
14
*
APB_DWIDTH
:
13
*
APB_DWIDTH
+
1
]
;
6
'h
20
:
CPWMl11
=
pwm_posedge_out_wire
[
15
*
APB_DWIDTH
:
14
*
APB_DWIDTH
+
1
]
;
6
'h
21
:
CPWMl11
=
pwm_negedge_out_wire
[
15
*
APB_DWIDTH
:
14
*
APB_DWIDTH
+
1
]
;
6
'h
24
:
CPWMl11
=
PWM_STRETCH
[
PWM_NUM
-
1
:
0
]
;
default
:
CPWMl11
=
0
;
endcase
end
end
endgenerate
generate
if
(
PWM_NUM
==
16
)
begin
:
CPWMIO1
always
@*
begin
case
(
PADDR
)
6
'h
02
:
CPWMl11
=
pwm_enable_out_wire
[
8
:
1
]
;
6
'h
03
:
CPWMl11
=
pwm_enable_out_wire
[
16
:
9
]
;
6
'h
04
:
CPWMl11
=
pwm_posedge_out_wire
[
1
*
APB_DWIDTH
:
0
*
APB_DWIDTH
+
1
]
;
6
'h
05
:
CPWMl11
=
pwm_negedge_out_wire
[
1
*
APB_DWIDTH
:
0
*
APB_DWIDTH
+
1
]
;
6
'h
06
:
CPWMl11
=
pwm_posedge_out_wire
[
2
*
APB_DWIDTH
:
1
*
APB_DWIDTH
+
1
]
;
6
'h
07
:
CPWMl11
=
pwm_negedge_out_wire
[
2
*
APB_DWIDTH
:
1
*
APB_DWIDTH
+
1
]
;
6
'h
08
:
CPWMl11
=
pwm_posedge_out_wire
[
3
*
APB_DWIDTH
:
2
*
APB_DWIDTH
+
1
]
;
6
'h
09
:
CPWMl11
=
pwm_negedge_out_wire
[
3
*
APB_DWIDTH
:
2
*
APB_DWIDTH
+
1
]
;
6
'h
0a
:
CPWMl11
=
pwm_posedge_out_wire
[
4
*
APB_DWIDTH
:
3
*
APB_DWIDTH
+
1
]
;
6
'h
0b
:
CPWMl11
=
pwm_negedge_out_wire
[
4
*
APB_DWIDTH
:
3
*
APB_DWIDTH
+
1
]
;
6
'h
0c
:
CPWMl11
=
pwm_posedge_out_wire
[
5
*
APB_DWIDTH
:
4
*
APB_DWIDTH
+
1
]
;
6
'h
0d
:
CPWMl11
=
pwm_negedge_out_wire
[
5
*
APB_DWIDTH
:
4
*
APB_DWIDTH
+
1
]
;
6
'h
0e
:
CPWMl11
=
pwm_posedge_out_wire
[
6
*
APB_DWIDTH
:
5
*
APB_DWIDTH
+
1
]
;
6
'h
0f
:
CPWMl11
=
pwm_negedge_out_wire
[
6
*
APB_DWIDTH
:
5
*
APB_DWIDTH
+
1
]
;
6
'h
10
:
CPWMl11
=
pwm_posedge_out_wire
[
7
*
APB_DWIDTH
:
6
*
APB_DWIDTH
+
1
]
;
6
'h
11
:
CPWMl11
=
pwm_negedge_out_wire
[
7
*
APB_DWIDTH
:
6
*
APB_DWIDTH
+
1
]
;
6
'h
12
:
CPWMl11
=
pwm_posedge_out_wire
[
8
*
APB_DWIDTH
:
7
*
APB_DWIDTH
+
1
]
;
6
'h
13
:
CPWMl11
=
pwm_negedge_out_wire
[
8
*
APB_DWIDTH
:
7
*
APB_DWIDTH
+
1
]
;
6
'h
14
:
CPWMl11
=
pwm_posedge_out_wire
[
9
*
APB_DWIDTH
:
8
*
APB_DWIDTH
+
1
]
;
6
'h
15
:
CPWMl11
=
pwm_negedge_out_wire
[
9
*
APB_DWIDTH
:
8
*
APB_DWIDTH
+
1
]
;
6
'h
16
:
CPWMl11
=
pwm_posedge_out_wire
[
10
*
APB_DWIDTH
:
9
*
APB_DWIDTH
+
1
]
;
6
'h
17
:
CPWMl11
=
pwm_negedge_out_wire
[
10
*
APB_DWIDTH
:
9
*
APB_DWIDTH
+
1
]
;
6
'h
18
:
CPWMl11
=
pwm_posedge_out_wire
[
11
*
APB_DWIDTH
:
10
*
APB_DWIDTH
+
1
]
;
6
'h
19
:
CPWMl11
=
pwm_negedge_out_wire
[
11
*
APB_DWIDTH
:
10
*
APB_DWIDTH
+
1
]
;
6
'h
1a
:
CPWMl11
=
pwm_posedge_out_wire
[
12
*
APB_DWIDTH
:
11
*
APB_DWIDTH
+
1
]
;
6
'h
1b
:
CPWMl11
=
pwm_negedge_out_wire
[
12
*
APB_DWIDTH
:
11
*
APB_DWIDTH
+
1
]
;
6
'h
1c
:
CPWMl11
=
pwm_posedge_out_wire
[
13
*
APB_DWIDTH
:
12
*
APB_DWIDTH
+
1
]
;
6
'h
1d
:
CPWMl11
=
pwm_negedge_out_wire
[
13
*
APB_DWIDTH
:
12
*
APB_DWIDTH
+
1
]
;
6
'h
1e
:
CPWMl11
=
pwm_posedge_out_wire
[
14
*
APB_DWIDTH
:
13
*
APB_DWIDTH
+
1
]
;
6
'h
1f
:
CPWMl11
=
pwm_negedge_out_wire
[
14
*
APB_DWIDTH
:
13
*
APB_DWIDTH
+
1
]
;
6
'h
20
:
CPWMl11
=
pwm_posedge_out_wire
[
15
*
APB_DWIDTH
:
14
*
APB_DWIDTH
+
1
]
;
6
'h
21
:
CPWMl11
=
pwm_negedge_out_wire
[
15
*
APB_DWIDTH
:
14
*
APB_DWIDTH
+
1
]
;
6
'h
22
:
CPWMl11
=
pwm_posedge_out_wire
[
16
*
APB_DWIDTH
:
15
*
APB_DWIDTH
+
1
]
;
6
'h
23
:
CPWMl11
=
pwm_negedge_out_wire
[
16
*
APB_DWIDTH
:
15
*
APB_DWIDTH
+
1
]
;
6
'h
24
:
CPWMl11
=
PWM_STRETCH
[
PWM_NUM
-
1
:
0
]
;
default
:
CPWMl11
=
0
;
endcase
end
end
endgenerate
generate
if
(
APB_DWIDTH
==
32
)
begin
assign
CPWMO0
=
(
PADDR
<=
1
)
?
CPWMI11
:
(
(
PADDR
==
57
)
?
{
31
'b
0
,
CPWMllOI
}
:
CPWMl11
)
;
end
else
if
(
APB_DWIDTH
==
16
)
begin
assign
CPWMO0
=
(
PADDR
<=
1
)
?
CPWMI11
:
(
(
PADDR
==
57
)
?
{
15
'b
0
,
CPWMllOI
}
:
CPWMl11
)
;
end
else
begin
assign
CPWMO0
=
(
PADDR
<=
1
)
?
CPWMI11
:
(
(
PADDR
==
57
)
?
{
7
'b
0
,
CPWMllOI
}
:
CPWMl11
)
;
end
endgenerate
endmodule
