// Actel Corporation Proprietary and Confidential
//  Copyright 2008 Actel Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE ACTEL LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
//  Revision Information:
// Jun09    Revision 4.1
// Aug10    Revision 4.2
// SVN Revision Information:
// SVN $Revision: 8508 $
// SVN $Date: 2009-06-15 16:49:49 -0700 (Mon, 15 Jun 2009) $
`timescale 1ns/1ns
module
CoreUARTapb_C0_CoreUARTapb_C0_0_Rx_async
(
CUARTII
,
CUARTIl
,
CUARTlI
,
CUARTII1
,
CUARTlI1
,
CUARTOl1
,
CUARTOOl
,
CUARTl0l
,
CUARTl01
,
CUARTO11
,
CUARTI11
,
CUARTI1l
,
CUARTllI
,
CUARTlOl
,
CUARTI0I
,
CUARTI01
,
CUARTO1l
,
CUARTIO0
,
CUARTI00
,
CUARTl00
)
;
parameter
SYNC_RESET
=
0
;
parameter
RX_FIFO
=
0
;
parameter
CUARTOIIl
=
0
;
parameter
CUARTIIIl
=
1
;
parameter
CUARTlIIl
=
2
;
parameter
CUARTOlIl
=
3
;
input
CUARTII
;
input
CUARTIl
;
input
CUARTlI
;
input
CUARTII1
;
input
CUARTlI1
;
input
CUARTOl1
;
input
CUARTOOl
;
input
CUARTl0l
;
input
CUARTO1l
;
input
CUARTl01
;
output
CUARTO11
;
output
CUARTI11
;
output
CUARTI1l
;
output
CUARTllI
;
output
[
7
:
0
]
CUARTlOl
;
output
CUARTI0I
;
output
CUARTI01
;
output
CUARTIO0
;
output
CUARTI00
;
output
CUARTl00
;
reg
CUARTI01
;
reg
CUARTI00
;
reg
CUARTO11
;
reg
CUARTI11
;
reg
CUARTI0I
;
wire
CUARTllI
;
reg
[
7
:
0
]
CUARTlOl
;
reg
[
1
:
0
]
CUARTll0
;
reg
[
3
:
0
]
CUARTIlIl
;
reg
CUARTllIl
;
reg
[
8
:
0
]
CUARTO0Il
;
reg
CUARTI0Il
;
reg
[
3
:
0
]
CUARTl0Il
;
reg
CUARTO1Il
;
reg
[
2
:
0
]
CUARTI1Il
;
reg
CUARTl1Il
;
reg
CUARTOOll
;
reg
CUARTI1l
;
reg
CUARTIO0
;
reg
[
3
:
0
]
CUARTIOll
;
wire
[
1
:
0
]
CUARTlOll
;
wire
[
1
:
0
]
CUARTOIll
;
wire
CUARTI1
;
wire
CUARTl1
;
assign
CUARTI1
=
(
SYNC_RESET
==
1
)
?
1
'b
1
:
CUARTlI
;
assign
CUARTl1
=
(
SYNC_RESET
==
1
)
?
CUARTlI
:
1
'b
1
;
always
@
(
posedge
CUARTII
or
negedge
CUARTI1
)
begin
:
CUARTIIll
if
(
(
!
CUARTI1
)
||
(
!
CUARTl1
)
)
begin
CUARTI1Il
<=
3
'b
111
;
end
else
begin
if
(
CUARTIl
==
1
'b
1
)
begin
CUARTI1Il
[
1
:
0
]
<=
CUARTI1Il
[
2
:
1
]
;
CUARTI1Il
[
2
]
<=
CUARTl01
;
end
end
end
always
@
(
CUARTI1Il
)
begin
case
(
CUARTI1Il
)
3
'b
000
:
begin
CUARTllIl
<=
1
'b
0
;
end
3
'b
001
:
begin
CUARTllIl
<=
1
'b
0
;
end
3
'b
010
:
begin
CUARTllIl
<=
1
'b
0
;
end
3
'b
011
:
begin
CUARTllIl
<=
1
'b
1
;
end
3
'b
100
:
begin
CUARTllIl
<=
1
'b
0
;
end
3
'b
101
:
begin
CUARTllIl
<=
1
'b
1
;
end
3
'b
110
:
begin
CUARTllIl
<=
1
'b
1
;
end
default
:
begin
CUARTllIl
<=
1
'b
1
;
end
endcase
end
always
@
(
posedge
CUARTII
or
negedge
CUARTI1
)
begin
:
CUARTlIll
if
(
(
!
CUARTI1
)
||
(
!
CUARTl1
)
)
begin
CUARTIlIl
<=
4
'b
0000
;
end
else
begin
if
(
CUARTIl
==
1
'b
1
)
begin
if
(
(
CUARTll0
==
CUARTOIIl
&
(
CUARTllIl
==
1
'b
1
|
CUARTIlIl
==
4
'b
1000
)
)
||
(
(
CUARTll0
==
CUARTOlIl
)
&&
(
CUARTIlIl
==
4
'b
0110
)
)
)
begin
CUARTIlIl
<=
4
'b
0000
;
end
else
begin
CUARTIlIl
<=
CUARTIlIl
+
1
'b
1
;
end
end
end
end
always
@
(
posedge
CUARTII
or
negedge
CUARTI1
)
begin
:
CUARTOlll
if
(
(
!
CUARTI1
)
||
(
!
CUARTl1
)
)
begin
CUARTO11
<=
1
'b
0
;
end
else
begin
if
(
CUARTIl
==
1
'b
1
)
begin
if
(
CUARTl1Il
==
1
'b
1
)
begin
CUARTO11
<=
1
'b
1
;
end
end
if
(
CUARTOOl
==
1
'b
1
)
begin
CUARTO11
<=
1
'b
0
;
end
end
end
always
@
(
posedge
CUARTII
or
negedge
CUARTI1
)
begin
:
CUARTIlll
if
(
(
!
CUARTI1
)
||
(
!
CUARTl1
)
)
begin
CUARTI01
<=
1
'b
0
;
end
else
if
(
CUARTIl
==
1
'b
1
)
begin
if
(
CUARTOOll
==
1
'b
1
)
begin
CUARTI01
<=
1
'b
1
;
end
else
if
(
CUARTO1l
==
1
'b
1
)
begin
CUARTI01
<=
1
'b
0
;
end
end
else
if
(
CUARTO1l
==
1
'b
1
)
begin
CUARTI01
<=
1
'b
0
;
end
else
begin
CUARTI01
<=
CUARTI01
;
end
end
always
@
(
posedge
CUARTII
or
negedge
CUARTI1
)
begin
if
(
(
!
CUARTI1
)
||
(
!
CUARTl1
)
)
begin
CUARTIOll
<=
4
'b
1001
;
end
else
begin
if
(
(
CUARTll0
==
CUARTOIIl
)
&&
(
CUARTIlIl
==
4
'b
1000
)
)
begin
case
(
{
CUARTII1
,
CUARTlI1
}
)
2
'b
00
:
CUARTIOll
<=
4
'b
0111
;
2
'b
01
:
CUARTIOll
<=
4
'b
1000
;
2
'b
10
:
CUARTIOll
<=
4
'b
1000
;
2
'b
11
:
CUARTIOll
<=
4
'b
1001
;
endcase
end
else
begin
CUARTIOll
<=
CUARTIOll
;
end
end
end
assign
CUARTl00
=
(
CUARTll0
==
CUARTOIIl
)
;
always
@
(
posedge
CUARTII
or
negedge
CUARTI1
)
begin
:
CUARTllll
if
(
(
!
CUARTI1
)
||
(
!
CUARTl1
)
)
begin
CUARTll0
<=
CUARTOIIl
;
CUARTlOl
<=
8
'b
00000000
;
CUARTl1Il
<=
1
'b
0
;
CUARTOOll
<=
1
'b
0
;
CUARTI00
<=
1
'b
0
;
end
else
begin
if
(
CUARTIl
==
1
'b
1
)
begin
CUARTl1Il
<=
1
'b
0
;
CUARTI00
<=
1
'b
0
;
CUARTOOll
<=
1
'b
0
;
case
(
CUARTll0
)
CUARTOIIl
:
begin
if
(
CUARTIlIl
==
4
'b
1000
)
begin
CUARTll0
<=
CUARTIIIl
;
end
else
begin
CUARTll0
<=
CUARTOIIl
;
end
end
CUARTIIIl
:
begin
if
(
CUARTl0Il
==
CUARTIOll
)
begin
CUARTll0
<=
CUARTlIIl
;
CUARTl1Il
<=
CUARTO1Il
;
if
(
CUARTO1Il
==
1
'b
0
)
begin
CUARTlOl
<=
{
(
CUARTII1
&
CUARTO0Il
[
7
]
)
,
CUARTO0Il
[
6
:
0
]
}
;
end
end
else
begin
CUARTll0
<=
CUARTIIIl
;
end
end
CUARTlIIl
:
begin
if
(
CUARTIlIl
==
4
'b
1110
)
begin
if
(
CUARTllIl
==
1
'b
0
)
begin
CUARTOOll
<=
1
'b
1
;
end
end
else
if
(
CUARTIlIl
==
4
'b
1111
)
begin
CUARTI00
<=
1
'b
1
;
CUARTll0
<=
CUARTOlIl
;
end
else
begin
CUARTll0
<=
CUARTlIIl
;
end
end
CUARTOlIl
:
begin
if
(
(
CUARTllIl
==
1
'b
1
)
||
(
CUARTIlIl
==
4
'b
0110
)
)
begin
CUARTll0
<=
CUARTOIIl
;
end
else
begin
CUARTll0
<=
CUARTOlIl
;
end
end
default
:
begin
CUARTll0
<=
CUARTOIIl
;
end
endcase
end
end
end
assign
CUARTlOll
=
{
CUARTII1
,
CUARTlI1
}
;
always
@
(
posedge
CUARTII
or
negedge
CUARTI1
)
begin
:
CUARTO0ll
if
(
(
!
CUARTI1
)
||
(
!
CUARTl1
)
)
begin
CUARTO0Il
[
8
:
0
]
<=
9
'b
000000000
;
CUARTl0Il
<=
4
'b
0000
;
end
else
begin
if
(
CUARTIl
==
1
'b
1
)
begin
if
(
CUARTll0
==
CUARTOIIl
)
begin
CUARTO0Il
[
8
:
0
]
<=
9
'b
000000000
;
CUARTl0Il
<=
4
'b
0000
;
end
else
if
(
CUARTIlIl
==
4
'b
1111
)
begin
CUARTl0Il
<=
CUARTl0Il
+
1
'b
1
;
case
(
CUARTlOll
)
2
'b
00
:
begin
CUARTO0Il
[
5
:
0
]
<=
CUARTO0Il
[
6
:
1
]
;
CUARTO0Il
[
6
]
<=
CUARTllIl
;
end
2
'b
11
:
begin
CUARTO0Il
[
7
:
0
]
<=
CUARTO0Il
[
8
:
1
]
;
CUARTO0Il
[
8
]
<=
CUARTllIl
;
end
default
:
begin
CUARTO0Il
[
6
:
0
]
<=
CUARTO0Il
[
7
:
1
]
;
CUARTO0Il
[
7
]
<=
CUARTllIl
;
end
endcase
end
end
end
end
always
@
(
posedge
CUARTII
or
negedge
CUARTI1
)
begin
:
CUARTI0ll
if
(
(
!
CUARTI1
)
||
(
!
CUARTl1
)
)
begin
CUARTI0Il
<=
1
'b
0
;
end
else
begin
if
(
CUARTIl
==
1
'b
1
)
begin
if
(
CUARTIlIl
==
4
'b
1111
&
CUARTlI1
==
1
'b
1
)
begin
CUARTI0Il
<=
CUARTI0Il
^
CUARTllIl
;
end
if
(
CUARTll0
==
CUARTlIIl
)
begin
CUARTI0Il
<=
1
'b
0
;
end
end
end
end
assign
CUARTOIll
=
{
CUARTII1
,
CUARTOl1
}
;
always
@
(
posedge
CUARTII
or
negedge
CUARTI1
)
begin
:
CUARTl0ll
if
(
(
!
CUARTI1
)
||
(
!
CUARTl1
)
)
begin
CUARTI11
<=
1
'b
0
;
end
else
begin
if
(
CUARTIl
==
1
'b
1
&
CUARTlI1
==
1
'b
1
&
CUARTIlIl
==
4
'b
1111
)
begin
case
(
CUARTOIll
)
2
'b
00
:
begin
if
(
CUARTl0Il
==
4
'b
0111
)
begin
CUARTI11
<=
CUARTI0Il
^
CUARTllIl
;
end
end
2
'b
01
:
begin
if
(
CUARTl0Il
==
4
'b
0111
)
begin
CUARTI11
<=
~
(
CUARTI0Il
^
CUARTllIl
)
;
end
end
2
'b
10
:
begin
if
(
CUARTl0Il
==
4
'b
1000
)
begin
CUARTI11
<=
CUARTI0Il
^
CUARTllIl
;
end
end
2
'b
11
:
begin
if
(
CUARTl0Il
==
4
'b
1000
)
begin
CUARTI11
<=
~
(
CUARTI0Il
^
CUARTllIl
)
;
end
end
default
:
begin
CUARTI11
<=
1
'b
0
;
end
endcase
end
if
(
CUARTl0l
==
1
'b
1
)
begin
CUARTI11
<=
1
'b
0
;
end
end
end
always
@
(
posedge
CUARTII
or
negedge
CUARTI1
)
begin
:
CUARTO1ll
if
(
(
!
CUARTI1
)
||
(
!
CUARTl1
)
)
begin
CUARTO1Il
<=
1
'b
0
;
CUARTI0I
<=
1
'b
1
;
CUARTI1l
<=
1
'b
0
;
CUARTIO0
<=
1
'b
0
;
end
else
begin
CUARTI0I
<=
1
'b
1
;
CUARTI1l
<=
1
'b
0
;
CUARTIO0
<=
1
'b
0
;
if
(
CUARTIl
==
1
'b
1
)
begin
if
(
CUARTII1
==
1
'b
1
)
begin
if
(
CUARTlI1
==
1
'b
1
)
begin
if
(
CUARTl0Il
==
4
'b
1001
&
CUARTll0
==
CUARTIIIl
)
begin
CUARTI0I
<=
1
'b
0
;
CUARTI1l
<=
1
'b
1
;
CUARTIO0
<=
1
'b
1
;
if
(
RX_FIFO
==
1
'b
0
)
begin
CUARTO1Il
<=
1
'b
1
;
end
end
end
else
begin
if
(
CUARTl0Il
==
4
'b
1000
&
CUARTll0
==
CUARTIIIl
)
begin
CUARTI0I
<=
1
'b
0
;
CUARTI1l
<=
1
'b
1
;
CUARTIO0
<=
1
'b
1
;
if
(
RX_FIFO
==
1
'b
0
)
begin
CUARTO1Il
<=
1
'b
1
;
end
end
end
end
else
begin
if
(
CUARTlI1
==
1
'b
1
)
begin
if
(
CUARTl0Il
==
4
'b
1000
&
CUARTll0
==
CUARTIIIl
)
begin
CUARTI0I
<=
1
'b
0
;
CUARTI1l
<=
1
'b
1
;
CUARTIO0
<=
1
'b
1
;
if
(
RX_FIFO
==
1
'b
0
)
begin
CUARTO1Il
<=
1
'b
1
;
end
end
end
else
begin
if
(
CUARTl0Il
==
4
'b
0111
&
CUARTll0
==
CUARTIIIl
)
begin
CUARTI0I
<=
1
'b
0
;
CUARTI1l
<=
1
'b
1
;
CUARTIO0
<=
1
'b
1
;
if
(
RX_FIFO
==
1
'b
0
)
begin
CUARTO1Il
<=
1
'b
1
;
end
end
end
end
end
if
(
CUARTOOl
==
1
'b
1
)
begin
CUARTO1Il
<=
1
'b
0
;
end
end
end
assign
CUARTllI
=
CUARTO1Il
;
endmodule
