//////////////////////////////////////////////////////////////////////
// Created by SmartDesign Tue Mar 12 08:59:57 2024
// Version: 2023.2 2023.2.0.10
//////////////////////////////////////////////////////////////////////

`timescale 1ns / 100ps

//////////////////////////////////////////////////////////////////////
// Component Description (Tcl) 
//////////////////////////////////////////////////////////////////////
/*
# Exporting Component Description of IO_C1 to TCL
# Family: SmartFusion2
# Part Number: M2S025-1VF256I
# Create and Configure the core component IO_C1
create_and_configure_core -core_vlnv {Actel:SgCore:IO:1.0.101} -component_name {IO_C1} -params {\
"DIFF_IOSTD_OK:false"  \
"IO_TYPE:INBUF"  \
"IOSTD:LVCMOS33"  \
"SINGLE_IOSTD_OK:true"  \
"VARIATION:SINGLE"  \
"WIDTH:1"   }
# Exporting Component Description of IO_C1 to TCL done
*/

// IO_C1
module IO_C1(
    // Inputs
    PAD_IN,
    // Outputs
    Y
);

//--------------------------------------------------------------------
// Input
//--------------------------------------------------------------------
input  [0:0] PAD_IN;
//--------------------------------------------------------------------
// Output
//--------------------------------------------------------------------
output [0:0] Y;
//--------------------------------------------------------------------
// Nets
//--------------------------------------------------------------------
wire   [0:0] PAD_IN;
wire   [0:0] Y_net_0;
wire   [0:0] Y_net_1;
//--------------------------------------------------------------------
// TiedOff Nets
//--------------------------------------------------------------------
wire         GND_net;
//--------------------------------------------------------------------
// Constant assignments
//--------------------------------------------------------------------
assign GND_net    = 1'b0;
//--------------------------------------------------------------------
// Top level output port assignments
//--------------------------------------------------------------------
assign Y_net_1[0] = Y_net_0[0];
assign Y[0:0]     = Y_net_1[0];
//--------------------------------------------------------------------
// Component instances
//--------------------------------------------------------------------
//--------IO_C1_IO_C1_0_IO   -   Actel:SgCore:IO:1.0.101
IO_C1_IO_C1_0_IO IO_C1_0(
        // Inputs
        .PAD_IN ( PAD_IN ),
        // Outputs
        .Y      ( Y_net_0 ) 
        );


endmodule
