// Actel Corporation Proprietary and Confidential
// Copyright 2013 Actel Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE ACTEL LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
// SVN Revision Information:
// SVN $Revision: 23120 $
// SVN $Date: 2014-07-17 15:26:23 +0100 (Thu, 17 Jul 2014) $
`timescale 1ns/1ps
module
CAHBLTIIlll
#
(
parameter
[
2
:
0
]
MEMSPACE
=
0
,
parameter
[
0
:
0
]
HADDR_SHG_CFG
=
1
,
parameter
[
15
:
0
]
CAHBLTI
=
0
,
parameter
[
16
:
0
]
CAHBLTIIO0
=
(
2
**
17
)
-
1
,
parameter
[
16
:
0
]
CAHBLTlIO0
=
(
2
**
17
)
-
1
,
parameter
[
16
:
0
]
CAHBLTlIlll
=
(
2
**
17
)
-
1
,
parameter
[
16
:
0
]
CAHBLTOllll
=
(
2
**
17
)
-
1
,
parameter
SYNC_RESET
=
0
)
(
input
HCLK,
input
HRESETN,
input
REMAP_M0,
input
[
31
:
0
]
HADDR_M0,
input
HMASTLOCK_M0,
input
[
2
:
0
]
HSIZE_M0,
input
HTRANS_M0,
input
HWRITE_M0,
input
[
31
:
0
]
HWDATA_M0,
output
wire
HRESP_M0,
output
wire
[
31
:
0
]
HRDATA_M0,
output
wire
HREADY_M0,
input
[
31
:
0
]
HADDR_M1,
input
HMASTLOCK_M1,
input
[
2
:
0
]
HSIZE_M1,
input
HTRANS_M1,
input
HWRITE_M1,
input
[
31
:
0
]
HWDATA_M1,
output
wire
HRESP_M1,
output
wire
[
31
:
0
]
HRDATA_M1,
output
wire
HREADY_M1,
input
[
31
:
0
]
HADDR_M2,
input
HMASTLOCK_M2,
input
[
2
:
0
]
HSIZE_M2,
input
HTRANS_M2,
input
HWRITE_M2,
input
[
31
:
0
]
HWDATA_M2,
output
wire
HRESP_M2,
output
wire
[
31
:
0
]
HRDATA_M2,
output
wire
HREADY_M2,
input
[
31
:
0
]
HADDR_M3,
input
HMASTLOCK_M3,
input
[
2
:
0
]
HSIZE_M3,
input
HTRANS_M3,
input
HWRITE_M3,
input
[
31
:
0
]
HWDATA_M3,
output
wire
HRESP_M3,
output
wire
[
31
:
0
]
HRDATA_M3,
output
wire
HREADY_M3,
input
[
31
:
0
]
HRDATA_S0,
input
HREADYOUT_S0,
input
HRESP_S0,
output
wire
HSEL_S0,
output
wire
[
31
:
0
]
HADDR_S0,
output
wire
[
2
:
0
]
HSIZE_S0,
output
wire
HTRANS_S0,
output
wire
HWRITE_S0,
output
wire
[
31
:
0
]
HWDATA_S0,
output
wire
HREADY_S0,
output
wire
HMASTLOCK_S0,
input
[
31
:
0
]
HRDATA_S1,
input
HREADYOUT_S1,
input
HRESP_S1,
output
wire
HSEL_S1,
output
wire
[
31
:
0
]
HADDR_S1,
output
wire
[
2
:
0
]
HSIZE_S1,
output
wire
HTRANS_S1,
output
wire
HWRITE_S1,
output
wire
[
31
:
0
]
HWDATA_S1,
output
wire
HREADY_S1,
output
wire
HMASTLOCK_S1,
input
[
31
:
0
]
HRDATA_S2,
input
HREADYOUT_S2,
input
HRESP_S2,
output
wire
HSEL_S2,
output
wire
[
31
:
0
]
HADDR_S2,
output
wire
[
2
:
0
]
HSIZE_S2,
output
wire
HTRANS_S2,
output
wire
HWRITE_S2,
output
wire
[
31
:
0
]
HWDATA_S2,
output
wire
HREADY_S2,
output
wire
HMASTLOCK_S2,
input
[
31
:
0
]
HRDATA_S3,
input
HREADYOUT_S3,
input
HRESP_S3,
output
wire
HSEL_S3,
output
wire
[
31
:
0
]
HADDR_S3,
output
wire
[
2
:
0
]
HSIZE_S3,
output
wire
HTRANS_S3,
output
wire
HWRITE_S3,
output
wire
[
31
:
0
]
HWDATA_S3,
output
wire
HREADY_S3,
output
wire
HMASTLOCK_S3,
input
[
31
:
0
]
HRDATA_S4,
input
HREADYOUT_S4,
input
HRESP_S4,
output
wire
HSEL_S4,
output
wire
[
31
:
0
]
HADDR_S4,
output
wire
[
2
:
0
]
HSIZE_S4,
output
wire
HTRANS_S4,
output
wire
HWRITE_S4,
output
wire
[
31
:
0
]
HWDATA_S4,
output
wire
HREADY_S4,
output
wire
HMASTLOCK_S4,
input
[
31
:
0
]
HRDATA_S5,
input
HREADYOUT_S5,
input
HRESP_S5,
output
wire
HSEL_S5,
output
wire
[
31
:
0
]
HADDR_S5,
output
wire
[
2
:
0
]
HSIZE_S5,
output
wire
HTRANS_S5,
output
wire
HWRITE_S5,
output
wire
[
31
:
0
]
HWDATA_S5,
output
wire
HREADY_S5,
output
wire
HMASTLOCK_S5,
input
[
31
:
0
]
HRDATA_S6,
input
HREADYOUT_S6,
input
HRESP_S6,
output
wire
HSEL_S6,
output
wire
[
31
:
0
]
HADDR_S6,
output
wire
[
2
:
0
]
HSIZE_S6,
output
wire
HTRANS_S6,
output
wire
HWRITE_S6,
output
wire
[
31
:
0
]
HWDATA_S6,
output
wire
HREADY_S6,
output
wire
HMASTLOCK_S6,
input
[
31
:
0
]
HRDATA_S7,
input
HREADYOUT_S7,
input
HRESP_S7,
output
wire
HSEL_S7,
output
wire
[
31
:
0
]
HADDR_S7,
output
wire
[
2
:
0
]
HSIZE_S7,
output
wire
HTRANS_S7,
output
wire
HWRITE_S7,
output
wire
[
31
:
0
]
HWDATA_S7,
output
wire
HREADY_S7,
output
wire
HMASTLOCK_S7,
input
[
31
:
0
]
HRDATA_S8,
input
HREADYOUT_S8,
input
HRESP_S8,
output
wire
HSEL_S8,
output
wire
[
31
:
0
]
HADDR_S8,
output
wire
[
2
:
0
]
HSIZE_S8,
output
wire
HTRANS_S8,
output
wire
HWRITE_S8,
output
wire
[
31
:
0
]
HWDATA_S8,
output
wire
HREADY_S8,
output
wire
HMASTLOCK_S8,
input
[
31
:
0
]
HRDATA_S9,
input
HREADYOUT_S9,
input
HRESP_S9,
output
wire
HSEL_S9,
output
wire
[
31
:
0
]
HADDR_S9,
output
wire
[
2
:
0
]
HSIZE_S9,
output
wire
HTRANS_S9,
output
wire
HWRITE_S9,
output
wire
[
31
:
0
]
HWDATA_S9,
output
wire
HREADY_S9,
output
wire
HMASTLOCK_S9,
input
[
31
:
0
]
HRDATA_S10,
input
HREADYOUT_S10,
input
HRESP_S10,
output
wire
HSEL_S10,
output
wire
[
31
:
0
]
HADDR_S10,
output
wire
[
2
:
0
]
HSIZE_S10,
output
wire
HTRANS_S10,
output
wire
HWRITE_S10,
output
wire
[
31
:
0
]
HWDATA_S10,
output
wire
HREADY_S10,
output
wire
HMASTLOCK_S10,
input
[
31
:
0
]
HRDATA_S11,
input
HREADYOUT_S11,
input
HRESP_S11,
output
wire
HSEL_S11,
output
wire
[
31
:
0
]
HADDR_S11,
output
wire
[
2
:
0
]
HSIZE_S11,
output
wire
HTRANS_S11,
output
wire
HWRITE_S11,
output
wire
[
31
:
0
]
HWDATA_S11,
output
wire
HREADY_S11,
output
wire
HMASTLOCK_S11,
input
[
31
:
0
]
HRDATA_S12,
input
HREADYOUT_S12,
input
HRESP_S12,
output
wire
HSEL_S12,
output
wire
[
31
:
0
]
HADDR_S12,
output
wire
[
2
:
0
]
HSIZE_S12,
output
wire
HTRANS_S12,
output
wire
HWRITE_S12,
output
wire
[
31
:
0
]
HWDATA_S12,
output
wire
HREADY_S12,
output
wire
HMASTLOCK_S12,
input
[
31
:
0
]
HRDATA_S13,
input
HREADYOUT_S13,
input
HRESP_S13,
output
wire
HSEL_S13,
output
wire
[
31
:
0
]
HADDR_S13,
output
wire
[
2
:
0
]
HSIZE_S13,
output
wire
HTRANS_S13,
output
wire
HWRITE_S13,
output
wire
[
31
:
0
]
HWDATA_S13,
output
wire
HREADY_S13,
output
wire
HMASTLOCK_S13,
input
[
31
:
0
]
HRDATA_S14,
input
HREADYOUT_S14,
input
HRESP_S14,
output
wire
HSEL_S14,
output
wire
[
31
:
0
]
HADDR_S14,
output
wire
[
2
:
0
]
HSIZE_S14,
output
wire
HTRANS_S14,
output
wire
HWRITE_S14,
output
wire
[
31
:
0
]
HWDATA_S14,
output
wire
HREADY_S14,
output
wire
HMASTLOCK_S14,
input
[
31
:
0
]
HRDATA_S15,
input
HREADYOUT_S15,
input
HRESP_S15,
output
wire
HSEL_S15,
output
wire
[
31
:
0
]
HADDR_S15,
output
wire
[
2
:
0
]
HSIZE_S15,
output
wire
HTRANS_S15,
output
wire
HWRITE_S15,
output
wire
[
31
:
0
]
HWDATA_S15,
output
wire
HREADY_S15,
output
wire
HMASTLOCK_S15,
input
[
31
:
0
]
HRDATA_S16,
input
HREADYOUT_S16,
input
HRESP_S16,
output
wire
HSEL_S16,
output
wire
[
31
:
0
]
HADDR_S16,
output
wire
[
2
:
0
]
HSIZE_S16,
output
wire
HTRANS_S16,
output
wire
HWRITE_S16,
output
wire
[
31
:
0
]
HWDATA_S16,
output
wire
HREADY_S16,
output
wire
HMASTLOCK_S16
)
;
wire
[
31
:
0
]
CAHBLTI11I
;
wire
CAHBLTlI0
;
wire
[
2
:
0
]
CAHBLTl11I
;
wire
CAHBLTOOOl
;
wire
CAHBLTIOOl
;
wire
CAHBLTOlO0
;
wire
CAHBLTIlO0
;
wire
CAHBLTllO0
;
wire
CAHBLTO0O0
;
wire
CAHBLTI0O0
;
wire
CAHBLTl0O0
;
wire
CAHBLTO1O0
;
wire
CAHBLTI1O0
;
wire
CAHBLTl1O0
;
wire
CAHBLTOOI0
;
wire
CAHBLTIOI0
;
wire
CAHBLTlOI0
;
wire
CAHBLTOII0
;
wire
CAHBLTIII0
;
wire
CAHBLTlII0
;
wire
CAHBLTOlI0
;
wire
CAHBLTIlI0
;
wire
CAHBLTllI0
;
wire
CAHBLTO0I0
;
wire
CAHBLTI0I0
;
wire
CAHBLTl0I0
;
wire
CAHBLTO1I0
;
wire
CAHBLTI1I0
;
wire
CAHBLTl1I0
;
wire
CAHBLTOOl0
;
wire
CAHBLTIOl0
;
wire
CAHBLTlOl0
;
wire
CAHBLTOIl0
;
wire
CAHBLTIIl0
;
wire
CAHBLTlIl0
;
wire
CAHBLTOll0
;
wire
CAHBLTIll0
;
wire
CAHBLTlll0
;
wire
CAHBLTO0l0
;
wire
CAHBLTI0l0
;
wire
CAHBLTl0l0
;
wire
CAHBLTO1l0
;
wire
CAHBLTI1l0
;
wire
CAHBLTl1l0
;
wire
CAHBLTOO00
;
wire
CAHBLTIO00
;
wire
CAHBLTlO00
;
wire
CAHBLTOI00
;
wire
CAHBLTII00
;
wire
CAHBLTlI00
;
wire
CAHBLTOl00
;
wire
CAHBLTIl00
;
wire
CAHBLTll00
;
wire
CAHBLTO000
;
wire
CAHBLTI000
;
wire
CAHBLTl000
;
wire
CAHBLTO100
;
wire
CAHBLTI100
;
wire
CAHBLTl100
;
wire
CAHBLTOO10
;
wire
CAHBLTIO10
;
wire
CAHBLTlO10
;
wire
CAHBLTOI10
;
wire
CAHBLTII10
;
wire
CAHBLTlI10
;
wire
CAHBLTOl10
;
wire
CAHBLTIl10
;
wire
CAHBLTll10
;
wire
CAHBLTO010
;
wire
CAHBLTI010
;
wire
CAHBLTl010
;
wire
CAHBLTO110
;
wire
CAHBLTI110
;
wire
CAHBLTl110
;
wire
CAHBLTOOO1
;
wire
CAHBLTIOO1
;
wire
CAHBLTlOO1
;
wire
CAHBLTOIO1
;
wire
CAHBLTIIO1
;
wire
CAHBLTlIO1
;
wire
CAHBLTOlO1
;
wire
CAHBLTIlO1
;
wire
CAHBLTllO1
;
wire
CAHBLTO0O1
;
wire
CAHBLTI0O1
;
wire
CAHBLTl0O1
;
wire
CAHBLTO1O1
;
wire
CAHBLTI1O1
;
wire
CAHBLTl1O1
;
wire
CAHBLTOOI1
;
wire
CAHBLTIOI1
;
wire
CAHBLTlOI1
;
wire
CAHBLTOII1
;
wire
CAHBLTIII1
;
wire
CAHBLTlII1
;
wire
CAHBLTOlI1
;
wire
CAHBLTIlI1
;
wire
CAHBLTllI1
;
wire
CAHBLTO0I1
;
wire
CAHBLTI0I1
;
wire
CAHBLTl0I1
;
wire
CAHBLTO1I1
;
wire
CAHBLTI1I1
;
wire
CAHBLTl1I1
;
wire
CAHBLTOOl1
;
wire
CAHBLTIOl1
;
wire
CAHBLTlOl1
;
wire
CAHBLTOIl1
;
wire
CAHBLTIIl1
;
wire
CAHBLTlIl1
;
wire
CAHBLTOll1
;
wire
CAHBLTIll1
;
wire
CAHBLTlll1
;
wire
CAHBLTO0l1
;
wire
CAHBLTI0l1
;
wire
CAHBLTl0l1
;
wire
CAHBLTO1l1
;
wire
CAHBLTI1l1
;
wire
CAHBLTl1l1
;
wire
CAHBLTOO01
;
wire
CAHBLTIO01
;
wire
CAHBLTlO01
;
wire
CAHBLTOI01
;
wire
CAHBLTII01
;
wire
CAHBLTlI01
;
wire
CAHBLTOl01
;
wire
CAHBLTIl01
;
wire
CAHBLTll01
;
wire
CAHBLTO001
;
wire
CAHBLTI001
;
wire
CAHBLTl001
;
wire
CAHBLTO101
;
wire
CAHBLTI101
;
wire
CAHBLTl101
;
wire
CAHBLTOO11
;
wire
CAHBLTIO11
;
wire
CAHBLTlO11
;
wire
CAHBLTOI11
;
wire
CAHBLTII11
;
wire
CAHBLTlI11
;
wire
CAHBLTOl11
;
wire
CAHBLTIl11
;
wire
CAHBLTll11
;
wire
CAHBLTO011
;
wire
CAHBLTI011
;
wire
CAHBLTl011
;
wire
CAHBLTO111
;
wire
CAHBLTI111
;
wire
CAHBLTl111
;
wire
CAHBLTOOOOI
;
wire
CAHBLTIOOOI
;
wire
CAHBLTlOOOI
;
wire
CAHBLTOIOOI
;
wire
CAHBLTIIOOI
;
wire
CAHBLTlIOOI
;
wire
CAHBLTOlOOI
;
wire
CAHBLTIlOOI
;
wire
CAHBLTllOOI
;
wire
CAHBLTO0OOI
;
wire
CAHBLTI0OOI
;
wire
CAHBLTl0OOI
;
wire
CAHBLTO1OOI
;
wire
CAHBLTI1OOI
;
wire
CAHBLTl1OOI
;
wire
CAHBLTOOIOI
;
wire
CAHBLTIOIOI
;
wire
CAHBLTlOIOI
;
wire
CAHBLTOIIOI
;
wire
CAHBLTIIIOI
;
wire
CAHBLTlIIOI
;
wire
CAHBLTOlIOI
;
wire
CAHBLTIlIOI
;
wire
CAHBLTllIOI
;
wire
CAHBLTO0IOI
;
wire
CAHBLTI0IOI
;
wire
CAHBLTl0IOI
;
wire
[
31
:
0
]
CAHBLTlOOl
;
wire
CAHBLTOl0
;
wire
[
2
:
0
]
CAHBLTOIOl
;
wire
CAHBLTIIOl
;
wire
CAHBLTlIOl
;
wire
CAHBLTO1IOI
;
wire
CAHBLTI1IOI
;
wire
CAHBLTl1IOI
;
wire
CAHBLTOOlOI
;
wire
CAHBLTIOlOI
;
wire
CAHBLTlOlOI
;
wire
CAHBLTOIlOI
;
wire
CAHBLTIIlOI
;
wire
CAHBLTlIlOI
;
wire
CAHBLTOllOI
;
wire
CAHBLTIllOI
;
wire
CAHBLTlllOI
;
wire
CAHBLTO0lOI
;
wire
CAHBLTI0lOI
;
wire
CAHBLTl0lOI
;
wire
CAHBLTO1lOI
;
wire
CAHBLTI1lOI
;
wire
CAHBLTl1lOI
;
wire
CAHBLTOO0OI
;
wire
CAHBLTIO0OI
;
wire
CAHBLTlO0OI
;
wire
CAHBLTOI0OI
;
wire
CAHBLTII0OI
;
wire
CAHBLTlI0OI
;
wire
CAHBLTOl0OI
;
wire
CAHBLTIl0OI
;
wire
CAHBLTll0OI
;
wire
CAHBLTO00OI
;
wire
CAHBLTI00OI
;
wire
CAHBLTl00OI
;
wire
CAHBLTO10OI
;
wire
CAHBLTI10OI
;
wire
CAHBLTl10OI
;
wire
CAHBLTOO1OI
;
wire
CAHBLTIO1OI
;
wire
CAHBLTlO1OI
;
wire
CAHBLTOI1OI
;
wire
CAHBLTII1OI
;
wire
CAHBLTlI1OI
;
wire
CAHBLTOl1OI
;
wire
CAHBLTIl1OI
;
wire
CAHBLTll1OI
;
wire
CAHBLTO01OI
;
wire
CAHBLTI01OI
;
wire
CAHBLTl01OI
;
wire
CAHBLTO11OI
;
wire
CAHBLTI11OI
;
wire
CAHBLTl11OI
;
wire
CAHBLTOOOII
;
wire
CAHBLTIOOII
;
wire
CAHBLTlOOII
;
wire
CAHBLTOIOII
;
wire
CAHBLTIIOII
;
wire
CAHBLTlIOII
;
wire
CAHBLTOlOII
;
wire
CAHBLTIlOII
;
wire
CAHBLTllOII
;
wire
CAHBLTO0OII
;
wire
CAHBLTI0OII
;
wire
CAHBLTl0OII
;
wire
CAHBLTO1OII
;
wire
CAHBLTI1OII
;
wire
CAHBLTl1OII
;
wire
CAHBLTOOIII
;
wire
CAHBLTIOIII
;
wire
CAHBLTlOIII
;
wire
CAHBLTOIIII
;
wire
CAHBLTIIIII
;
wire
CAHBLTlIIII
;
wire
CAHBLTOlIII
;
wire
CAHBLTIlIII
;
wire
CAHBLTllIII
;
wire
CAHBLTO0III
;
wire
CAHBLTI0III
;
wire
CAHBLTl0III
;
wire
CAHBLTO1III
;
wire
CAHBLTI1III
;
wire
CAHBLTl1III
;
wire
CAHBLTOOlII
;
wire
CAHBLTIOlII
;
wire
CAHBLTlOlII
;
wire
CAHBLTOIlII
;
wire
CAHBLTIIlII
;
wire
CAHBLTlIlII
;
wire
CAHBLTOllII
;
wire
CAHBLTIllII
;
wire
CAHBLTlllII
;
wire
CAHBLTO0lII
;
wire
CAHBLTI0lII
;
wire
CAHBLTl0lII
;
wire
CAHBLTO1lII
;
wire
CAHBLTI1lII
;
wire
CAHBLTl1lII
;
wire
CAHBLTOO0II
;
wire
CAHBLTIO0II
;
wire
CAHBLTlO0II
;
wire
CAHBLTOI0II
;
wire
CAHBLTII0II
;
wire
CAHBLTlI0II
;
wire
CAHBLTOl0II
;
wire
CAHBLTIl0II
;
wire
CAHBLTll0II
;
wire
CAHBLTO00II
;
wire
CAHBLTI00II
;
wire
CAHBLTl00II
;
wire
CAHBLTO10II
;
wire
CAHBLTI10II
;
wire
CAHBLTl10II
;
wire
CAHBLTOO1II
;
wire
CAHBLTIO1II
;
wire
CAHBLTlO1II
;
wire
CAHBLTOI1II
;
wire
CAHBLTII1II
;
wire
CAHBLTlI1II
;
wire
CAHBLTOl1II
;
wire
CAHBLTIl1II
;
wire
CAHBLTll1II
;
wire
CAHBLTO01II
;
wire
CAHBLTI01II
;
wire
CAHBLTl01II
;
wire
CAHBLTO11II
;
wire
CAHBLTI11II
;
wire
CAHBLTl11II
;
wire
CAHBLTOOOlI
;
wire
CAHBLTIOOlI
;
wire
CAHBLTlOOlI
;
wire
CAHBLTOIOlI
;
wire
CAHBLTIIOlI
;
wire
CAHBLTlIOlI
;
wire
CAHBLTOlOlI
;
wire
CAHBLTIlOlI
;
wire
CAHBLTllOlI
;
wire
CAHBLTO0OlI
;
wire
CAHBLTI0OlI
;
wire
CAHBLTl0OlI
;
wire
CAHBLTO1OlI
;
wire
CAHBLTI1OlI
;
wire
CAHBLTl1OlI
;
wire
CAHBLTOOIlI
;
wire
CAHBLTIOIlI
;
wire
CAHBLTlOIlI
;
wire
CAHBLTOIIlI
;
wire
CAHBLTIIIlI
;
wire
CAHBLTlIIlI
;
wire
CAHBLTOlIlI
;
wire
CAHBLTIlIlI
;
wire
CAHBLTllIlI
;
wire
CAHBLTO0IlI
;
wire
CAHBLTI0IlI
;
wire
CAHBLTl0IlI
;
wire
CAHBLTO1IlI
;
wire
CAHBLTI1IlI
;
wire
CAHBLTl1IlI
;
wire
CAHBLTOOllI
;
wire
CAHBLTIOllI
;
wire
CAHBLTlOllI
;
wire
CAHBLTOIllI
;
wire
CAHBLTIIllI
;
wire
CAHBLTlIllI
;
wire
CAHBLTOlllI
;
wire
CAHBLTIlllI
;
wire
CAHBLTllllI
;
wire
CAHBLTO0llI
;
wire
CAHBLTI0llI
;
wire
CAHBLTl0llI
;
wire
CAHBLTO1llI
;
wire
CAHBLTI1llI
;
wire
CAHBLTl1llI
;
wire
CAHBLTOO0lI
;
wire
CAHBLTIO0lI
;
wire
CAHBLTlO0lI
;
wire
[
31
:
0
]
CAHBLTOlOl
;
wire
CAHBLTIl0
;
wire
[
2
:
0
]
CAHBLTIlOl
;
wire
CAHBLTllOl
;
wire
CAHBLTO0Ol
;
wire
CAHBLTIllll
;
wire
CAHBLTlllll
;
wire
CAHBLTO0lll
;
wire
CAHBLTI0lll
;
wire
CAHBLTl0lll
;
wire
CAHBLTO1lll
;
wire
CAHBLTI1lll
;
wire
CAHBLTl1lll
;
wire
CAHBLTOO0ll
;
wire
CAHBLTIO0ll
;
wire
CAHBLTlO0ll
;
wire
CAHBLTOI0ll
;
wire
CAHBLTII0ll
;
wire
CAHBLTlI0ll
;
wire
CAHBLTOl0ll
;
wire
CAHBLTIl0ll
;
wire
CAHBLTll0ll
;
wire
CAHBLTO00ll
;
wire
CAHBLTI00ll
;
wire
CAHBLTl00ll
;
wire
CAHBLTO10ll
;
wire
CAHBLTI10ll
;
wire
CAHBLTl10ll
;
wire
CAHBLTOO1ll
;
wire
CAHBLTIO1ll
;
wire
CAHBLTlO1ll
;
wire
CAHBLTOI1ll
;
wire
CAHBLTII1ll
;
wire
CAHBLTlI1ll
;
wire
CAHBLTOl1ll
;
wire
CAHBLTIl1ll
;
wire
CAHBLTll1ll
;
wire
CAHBLTO01ll
;
wire
CAHBLTI01ll
;
wire
CAHBLTl01ll
;
wire
CAHBLTO11ll
;
wire
CAHBLTI11ll
;
wire
CAHBLTl11ll
;
wire
CAHBLTOOO0l
;
wire
CAHBLTIOO0l
;
wire
CAHBLTlOO0l
;
wire
CAHBLTOIO0l
;
wire
CAHBLTIIO0l
;
wire
CAHBLTlIO0l
;
wire
CAHBLTOlO0l
;
wire
CAHBLTIlO0l
;
wire
CAHBLTllO0l
;
wire
CAHBLTO0O0l
;
wire
CAHBLTI0O0l
;
wire
CAHBLTl0O0l
;
wire
CAHBLTO1O0l
;
wire
CAHBLTI1O0l
;
wire
CAHBLTl1O0l
;
wire
CAHBLTOOI0l
;
wire
CAHBLTIOI0l
;
wire
CAHBLTlOI0l
;
wire
CAHBLTOII0l
;
wire
CAHBLTIII0l
;
wire
CAHBLTlII0l
;
wire
CAHBLTOlI0l
;
wire
CAHBLTIlI0l
;
wire
CAHBLTllI0l
;
wire
CAHBLTO0I0l
;
wire
CAHBLTI0I0l
;
wire
CAHBLTl0I0l
;
wire
CAHBLTO1I0l
;
wire
CAHBLTI1I0l
;
wire
CAHBLTl1I0l
;
wire
CAHBLTOOl0l
;
wire
CAHBLTIOl0l
;
wire
CAHBLTlOl0l
;
wire
CAHBLTOIl0l
;
wire
CAHBLTIIl0l
;
wire
CAHBLTlIl0l
;
wire
CAHBLTOll0l
;
wire
CAHBLTIll0l
;
wire
CAHBLTlll0l
;
wire
CAHBLTO0l0l
;
wire
CAHBLTI0l0l
;
wire
CAHBLTl0l0l
;
wire
CAHBLTO1l0l
;
wire
CAHBLTI1l0l
;
wire
CAHBLTl1l0l
;
wire
CAHBLTOO00l
;
wire
CAHBLTIO00l
;
wire
CAHBLTlO00l
;
wire
CAHBLTOI00l
;
wire
CAHBLTII00l
;
wire
CAHBLTlI00l
;
wire
CAHBLTOl00l
;
wire
CAHBLTIl00l
;
wire
CAHBLTll00l
;
wire
CAHBLTO000l
;
wire
CAHBLTI000l
;
wire
CAHBLTl000l
;
wire
CAHBLTO100l
;
wire
CAHBLTI100l
;
wire
CAHBLTl100l
;
wire
CAHBLTOO10l
;
wire
CAHBLTIO10l
;
wire
CAHBLTlO10l
;
wire
CAHBLTOI10l
;
wire
CAHBLTII10l
;
wire
CAHBLTlI10l
;
wire
CAHBLTOl10l
;
wire
CAHBLTIl10l
;
wire
CAHBLTll10l
;
wire
CAHBLTO010l
;
wire
CAHBLTI010l
;
wire
CAHBLTl010l
;
wire
CAHBLTO110l
;
wire
CAHBLTI110l
;
wire
CAHBLTl110l
;
wire
CAHBLTOOO1l
;
wire
CAHBLTIOO1l
;
wire
CAHBLTlOO1l
;
wire
CAHBLTOIO1l
;
wire
CAHBLTIIO1l
;
wire
CAHBLTlIO1l
;
wire
CAHBLTOlO1l
;
wire
CAHBLTIlO1l
;
wire
CAHBLTllO1l
;
wire
CAHBLTO0O1l
;
wire
CAHBLTI0O1l
;
wire
CAHBLTl0O1l
;
wire
CAHBLTO1O1l
;
wire
CAHBLTI1O1l
;
wire
CAHBLTl1O1l
;
wire
CAHBLTOOI1l
;
wire
CAHBLTIOI1l
;
wire
CAHBLTlOI1l
;
wire
CAHBLTOII1l
;
wire
CAHBLTIII1l
;
wire
CAHBLTlII1l
;
wire
CAHBLTOlI1l
;
wire
CAHBLTIlI1l
;
wire
CAHBLTllI1l
;
wire
CAHBLTO0I1l
;
wire
CAHBLTI0I1l
;
wire
CAHBLTl0I1l
;
wire
CAHBLTO1I1l
;
wire
CAHBLTI1I1l
;
wire
CAHBLTl1I1l
;
wire
CAHBLTOOl1l
;
wire
CAHBLTIOl1l
;
wire
CAHBLTlOl1l
;
wire
CAHBLTOIl1l
;
wire
CAHBLTIIl1l
;
wire
CAHBLTlIl1l
;
wire
CAHBLTOll1l
;
wire
CAHBLTIll1l
;
wire
CAHBLTlll1l
;
wire
CAHBLTO0l1l
;
wire
CAHBLTI0l1l
;
wire
CAHBLTl0l1l
;
wire
CAHBLTO1l1l
;
wire
CAHBLTI1l1l
;
wire
CAHBLTl1l1l
;
wire
CAHBLTOO01l
;
wire
CAHBLTIO01l
;
wire
CAHBLTlO01l
;
wire
CAHBLTOI01l
;
wire
CAHBLTII01l
;
wire
CAHBLTlI01l
;
wire
CAHBLTOl01l
;
wire
CAHBLTIl01l
;
wire
CAHBLTll01l
;
wire
CAHBLTO001l
;
wire
CAHBLTI001l
;
wire
CAHBLTl001l
;
wire
CAHBLTO101l
;
wire
[
31
:
0
]
CAHBLTI0Ol
;
wire
CAHBLTll0
;
wire
[
2
:
0
]
CAHBLTl0Ol
;
wire
CAHBLTO1Ol
;
wire
CAHBLTI1Ol
;
wire
CAHBLTI101l
;
wire
CAHBLTl101l
;
wire
CAHBLTOO11l
;
wire
CAHBLTIO11l
;
wire
CAHBLTlO11l
;
wire
CAHBLTOI11l
;
wire
CAHBLTII11l
;
wire
CAHBLTlI11l
;
wire
CAHBLTOl11l
;
wire
CAHBLTIl11l
;
wire
CAHBLTll11l
;
wire
CAHBLTO011l
;
wire
CAHBLTI011l
;
wire
CAHBLTl011l
;
wire
CAHBLTO111l
;
wire
CAHBLTI111l
;
wire
CAHBLTl111l
;
wire
CAHBLTOOOO0
;
wire
CAHBLTIOOO0
;
wire
CAHBLTlOOO0
;
wire
CAHBLTOIOO0
;
wire
CAHBLTIIOO0
;
wire
CAHBLTlIOO0
;
wire
CAHBLTOlOO0
;
wire
CAHBLTIlOO0
;
wire
CAHBLTllOO0
;
wire
CAHBLTO0OO0
;
wire
CAHBLTI0OO0
;
wire
CAHBLTl0OO0
;
wire
CAHBLTO1OO0
;
wire
CAHBLTI1OO0
;
wire
CAHBLTl1OO0
;
wire
CAHBLTOOIO0
;
wire
CAHBLTIOIO0
;
wire
CAHBLTlOIO0
;
wire
CAHBLTOIIO0
;
wire
CAHBLTIIIO0
;
wire
CAHBLTlIIO0
;
wire
CAHBLTOlIO0
;
wire
CAHBLTIlIO0
;
wire
CAHBLTllIO0
;
wire
CAHBLTO0IO0
;
wire
CAHBLTI0IO0
;
wire
CAHBLTl0IO0
;
wire
CAHBLTO1IO0
;
wire
CAHBLTI1IO0
;
wire
CAHBLTl1IO0
;
wire
CAHBLTOOlO0
;
wire
CAHBLTIOlO0
;
wire
CAHBLTlOlO0
;
wire
CAHBLTOIlO0
;
wire
CAHBLTIIlO0
;
wire
CAHBLTlIlO0
;
wire
CAHBLTOllO0
;
wire
CAHBLTIllO0
;
wire
CAHBLTlllO0
;
wire
CAHBLTO0lO0
;
wire
CAHBLTI0lO0
;
wire
CAHBLTl0lO0
;
wire
CAHBLTO1lO0
;
wire
CAHBLTI1lO0
;
wire
CAHBLTl1lO0
;
wire
CAHBLTOO0O0
;
wire
CAHBLTIO0O0
;
wire
CAHBLTlO0O0
;
wire
CAHBLTOI0O0
;
wire
CAHBLTII0O0
;
wire
CAHBLTlI0O0
;
wire
CAHBLTOl0O0
;
wire
CAHBLTIl0O0
;
wire
CAHBLTll0O0
;
wire
CAHBLTO00O0
;
wire
CAHBLTI00O0
;
wire
CAHBLTl00O0
;
wire
CAHBLTO10O0
;
wire
CAHBLTI10O0
;
wire
CAHBLTl10O0
;
wire
CAHBLTOO1O0
;
wire
CAHBLTIO1O0
;
wire
CAHBLTlO1O0
;
wire
CAHBLTOI1O0
;
wire
CAHBLTII1O0
;
wire
CAHBLTlI1O0
;
wire
CAHBLTOl1O0
;
wire
CAHBLTIl1O0
;
wire
CAHBLTll1O0
;
wire
CAHBLTO01O0
;
wire
CAHBLTI01O0
;
wire
CAHBLTl01O0
;
wire
CAHBLTO11O0
;
wire
CAHBLTI11O0
;
wire
CAHBLTl11O0
;
wire
CAHBLTOOOI0
;
wire
CAHBLTIOOI0
;
wire
CAHBLTlOOI0
;
wire
CAHBLTOIOI0
;
wire
CAHBLTIIOI0
;
wire
CAHBLTlIOI0
;
wire
CAHBLTOlOI0
;
wire
CAHBLTIlOI0
;
wire
CAHBLTllOI0
;
wire
CAHBLTO0OI0
;
wire
CAHBLTI0OI0
;
wire
CAHBLTl0OI0
;
wire
CAHBLTO1OI0
;
wire
CAHBLTI1OI0
;
wire
CAHBLTl1OI0
;
wire
CAHBLTOOII0
;
wire
CAHBLTIOII0
;
wire
CAHBLTlOII0
;
wire
CAHBLTOIII0
;
wire
CAHBLTIIII0
;
wire
CAHBLTlIII0
;
wire
CAHBLTOlII0
;
wire
CAHBLTIlII0
;
wire
CAHBLTllII0
;
wire
CAHBLTO0II0
;
wire
CAHBLTI0II0
;
wire
CAHBLTl0II0
;
wire
CAHBLTO1II0
;
wire
CAHBLTI1II0
;
wire
CAHBLTl1II0
;
wire
CAHBLTOOlI0
;
wire
CAHBLTIOlI0
;
wire
CAHBLTlOlI0
;
wire
CAHBLTOIlI0
;
wire
CAHBLTIIlI0
;
wire
CAHBLTlIlI0
;
wire
CAHBLTOllI0
;
wire
CAHBLTIllI0
;
wire
CAHBLTlllI0
;
wire
CAHBLTO0lI0
;
wire
CAHBLTI0lI0
;
wire
CAHBLTl0lI0
;
wire
CAHBLTO1lI0
;
wire
CAHBLTI1lI0
;
wire
CAHBLTl1lI0
;
wire
CAHBLTOO0I0
;
wire
CAHBLTIO0I0
;
wire
CAHBLTlO0I0
;
wire
CAHBLTOI0I0
;
wire
CAHBLTII0I0
;
wire
CAHBLTlI0I0
;
wire
CAHBLTOl0I0
;
wire
CAHBLTIl0I0
;
wire
CAHBLTll0I0
;
wire
CAHBLTO00I0
;
wire
CAHBLTI00I0
;
wire
CAHBLTl00I0
;
wire
CAHBLTO10I0
;
wire
CAHBLTI10I0
;
wire
CAHBLTl10I0
;
wire
CAHBLTOO1I0
;
wire
CAHBLTIO1I0
;
wire
CAHBLTlO1I0
;
wire
CAHBLTOI1I0
;
wire
CAHBLTII1I0
;
wire
CAHBLTlI1I0
;
wire
CAHBLTOl1I0
;
wire
CAHBLTIl1I0
;
wire
CAHBLTll1I0
;
wire
CAHBLTO01I0
;
wire
CAHBLTI01I0
;
wire
CAHBLTl01I0
;
wire
CAHBLTO11I0
;
wire
CAHBLTI11I0
;
wire
CAHBLTl11I0
;
wire
CAHBLTOOOl0
;
wire
CAHBLTIOOl0
;
wire
CAHBLTlOOl0
;
wire
CAHBLTOIOl0
;
wire
[
31
:
0
]
CAHBLTOI0lI
;
wire
[
31
:
0
]
CAHBLTII0lI
;
wire
[
31
:
0
]
CAHBLTlI0lI
;
wire
[
31
:
0
]
CAHBLTOl0lI
;
wire
[
31
:
0
]
CAHBLTIl0lI
;
wire
[
31
:
0
]
CAHBLTll0lI
;
wire
[
31
:
0
]
CAHBLTO00lI
;
wire
[
31
:
0
]
CAHBLTI00lI
;
wire
[
31
:
0
]
CAHBLTl00lI
;
wire
[
31
:
0
]
CAHBLTO10lI
;
wire
[
31
:
0
]
CAHBLTI10lI
;
wire
[
31
:
0
]
CAHBLTl10lI
;
wire
[
31
:
0
]
CAHBLTOO1lI
;
wire
[
31
:
0
]
CAHBLTIO1lI
;
wire
[
31
:
0
]
CAHBLTlO1lI
;
wire
[
31
:
0
]
CAHBLTOI1lI
;
wire
[
31
:
0
]
CAHBLTII1lI
;
wire
[
31
:
0
]
CAHBLTlI1lI
;
wire
[
31
:
0
]
CAHBLTOl1lI
;
wire
[
31
:
0
]
CAHBLTIl1lI
;
wire
[
31
:
0
]
CAHBLTll1lI
;
wire
[
31
:
0
]
CAHBLTO01lI
;
wire
[
31
:
0
]
CAHBLTI01lI
;
wire
[
31
:
0
]
CAHBLTl01lI
;
wire
[
31
:
0
]
CAHBLTO11lI
;
wire
[
31
:
0
]
CAHBLTI11lI
;
wire
[
31
:
0
]
CAHBLTl11lI
;
wire
[
31
:
0
]
CAHBLTOOO0I
;
wire
[
31
:
0
]
CAHBLTIOO0I
;
wire
[
31
:
0
]
CAHBLTlOO0I
;
wire
[
31
:
0
]
CAHBLTOIO0I
;
wire
[
31
:
0
]
CAHBLTIIO0I
;
wire
[
31
:
0
]
CAHBLTlIO0I
;
wire
[
31
:
0
]
CAHBLTOlO0I
;
wire
[
31
:
0
]
CAHBLTIIOl0
;
wire
[
31
:
0
]
CAHBLTlIOl0
;
wire
[
31
:
0
]
CAHBLTOlOl0
;
wire
[
31
:
0
]
CAHBLTIlOl0
;
wire
[
31
:
0
]
CAHBLTllOl0
;
wire
[
31
:
0
]
CAHBLTO0Ol0
;
wire
[
31
:
0
]
CAHBLTI0Ol0
;
wire
[
31
:
0
]
CAHBLTl0Ol0
;
wire
[
31
:
0
]
CAHBLTO1Ol0
;
wire
[
31
:
0
]
CAHBLTI1Ol0
;
wire
[
31
:
0
]
CAHBLTl1Ol0
;
wire
[
31
:
0
]
CAHBLTOOIl0
;
wire
[
31
:
0
]
CAHBLTIOIl0
;
wire
[
31
:
0
]
CAHBLTlOIl0
;
wire
[
31
:
0
]
CAHBLTOIIl0
;
wire
[
31
:
0
]
CAHBLTIIIl0
;
wire
[
31
:
0
]
CAHBLTlIIl0
;
wire
[
31
:
0
]
CAHBLTOlIl0
;
wire
[
31
:
0
]
CAHBLTIlIl0
;
wire
[
31
:
0
]
CAHBLTllIl0
;
wire
[
31
:
0
]
CAHBLTO0Il0
;
wire
[
31
:
0
]
CAHBLTI0Il0
;
wire
[
31
:
0
]
CAHBLTl0Il0
;
wire
[
31
:
0
]
CAHBLTO1Il0
;
wire
[
31
:
0
]
CAHBLTI1Il0
;
wire
[
31
:
0
]
CAHBLTl1Il0
;
wire
[
31
:
0
]
CAHBLTOOll0
;
wire
[
31
:
0
]
CAHBLTIOll0
;
wire
[
31
:
0
]
CAHBLTlOll0
;
wire
[
31
:
0
]
CAHBLTOIll0
;
wire
[
31
:
0
]
CAHBLTIIll0
;
wire
[
31
:
0
]
CAHBLTlIll0
;
wire
[
31
:
0
]
CAHBLTOlll0
;
wire
[
31
:
0
]
CAHBLTIlll0
;
wire
CAHBLTIlO0I
;
wire
CAHBLTllO0I
;
wire
CAHBLTO0O0I
;
wire
CAHBLTI0O0I
;
wire
CAHBLTl0O0I
;
wire
CAHBLTO1O0I
;
wire
CAHBLTI1O0I
;
wire
CAHBLTl1O0I
;
wire
CAHBLTOOI0I
;
wire
CAHBLTIOI0I
;
wire
CAHBLTlOI0I
;
wire
CAHBLTOII0I
;
wire
CAHBLTIII0I
;
wire
CAHBLTlII0I
;
wire
CAHBLTOlI0I
;
wire
CAHBLTIlI0I
;
wire
CAHBLTllI0I
;
wire
CAHBLTO0I0I
;
wire
CAHBLTI0I0I
;
wire
CAHBLTl0I0I
;
wire
CAHBLTO1I0I
;
wire
CAHBLTI1I0I
;
wire
CAHBLTl1I0I
;
wire
CAHBLTOOl0I
;
wire
CAHBLTIOl0I
;
wire
CAHBLTlOl0I
;
wire
CAHBLTOIl0I
;
wire
CAHBLTIIl0I
;
wire
CAHBLTlIl0I
;
wire
CAHBLTOll0I
;
wire
CAHBLTIll0I
;
wire
CAHBLTlll0I
;
wire
CAHBLTO0l0I
;
wire
CAHBLTI0l0I
;
wire
CAHBLTllll0
;
wire
CAHBLTO0ll0
;
wire
CAHBLTI0ll0
;
wire
CAHBLTl0ll0
;
wire
CAHBLTO1ll0
;
wire
CAHBLTI1ll0
;
wire
CAHBLTl1ll0
;
wire
CAHBLTOO0l0
;
wire
CAHBLTIO0l0
;
wire
CAHBLTlO0l0
;
wire
CAHBLTOI0l0
;
wire
CAHBLTII0l0
;
wire
CAHBLTlI0l0
;
wire
CAHBLTOl0l0
;
wire
CAHBLTIl0l0
;
wire
CAHBLTll0l0
;
wire
CAHBLTO00l0
;
wire
CAHBLTI00l0
;
wire
CAHBLTl00l0
;
wire
CAHBLTO10l0
;
wire
CAHBLTI10l0
;
wire
CAHBLTl10l0
;
wire
CAHBLTOO1l0
;
wire
CAHBLTIO1l0
;
wire
CAHBLTlO1l0
;
wire
CAHBLTOI1l0
;
wire
CAHBLTII1l0
;
wire
CAHBLTlI1l0
;
wire
CAHBLTOl1l0
;
wire
CAHBLTIl1l0
;
wire
CAHBLTll1l0
;
wire
CAHBLTO01l0
;
wire
CAHBLTI01l0
;
wire
CAHBLTl01l0
;
wire
CAHBLTl0l0I
;
wire
CAHBLTO1l0I
;
wire
CAHBLTI1l0I
;
wire
CAHBLTl1l0I
;
wire
CAHBLTOO00I
;
wire
CAHBLTIO00I
;
wire
CAHBLTlO00I
;
wire
CAHBLTOI00I
;
wire
CAHBLTII00I
;
wire
CAHBLTlI00I
;
wire
CAHBLTOl00I
;
wire
CAHBLTIl00I
;
wire
CAHBLTll00I
;
wire
CAHBLTO000I
;
wire
CAHBLTI000I
;
wire
CAHBLTl000I
;
wire
CAHBLTO100I
;
wire
CAHBLTI100I
;
wire
CAHBLTl100I
;
wire
CAHBLTOO10I
;
wire
CAHBLTIO10I
;
wire
CAHBLTlO10I
;
wire
CAHBLTOI10I
;
wire
CAHBLTII10I
;
wire
CAHBLTlI10I
;
wire
CAHBLTOl10I
;
wire
CAHBLTIl10I
;
wire
CAHBLTll10I
;
wire
CAHBLTO010I
;
wire
CAHBLTI010I
;
wire
CAHBLTl010I
;
wire
CAHBLTO110I
;
wire
CAHBLTI110I
;
wire
CAHBLTl110I
;
wire
[
31
:
0
]
CAHBLTOOO1I
;
wire
[
31
:
0
]
CAHBLTIOO1I
;
wire
[
31
:
0
]
CAHBLTlOO1I
;
wire
[
31
:
0
]
CAHBLTOIO1I
;
wire
[
31
:
0
]
CAHBLTIIO1I
;
wire
[
31
:
0
]
CAHBLTlIO1I
;
wire
[
31
:
0
]
CAHBLTOlO1I
;
wire
[
31
:
0
]
CAHBLTIlO1I
;
wire
[
31
:
0
]
CAHBLTllO1I
;
wire
[
31
:
0
]
CAHBLTO0O1I
;
wire
[
31
:
0
]
CAHBLTI0O1I
;
wire
[
31
:
0
]
CAHBLTl0O1I
;
wire
[
31
:
0
]
CAHBLTO1O1I
;
wire
[
31
:
0
]
CAHBLTI1O1I
;
wire
[
31
:
0
]
CAHBLTl1O1I
;
wire
[
31
:
0
]
CAHBLTOOI1I
;
wire
[
31
:
0
]
CAHBLTIOI1I
;
wire
[
31
:
0
]
CAHBLTlOI1I
;
wire
[
31
:
0
]
CAHBLTOII1I
;
wire
[
31
:
0
]
CAHBLTIII1I
;
wire
[
31
:
0
]
CAHBLTlII1I
;
wire
[
31
:
0
]
CAHBLTOlI1I
;
wire
[
31
:
0
]
CAHBLTIlI1I
;
wire
[
31
:
0
]
CAHBLTllI1I
;
wire
[
31
:
0
]
CAHBLTO0I1I
;
wire
[
31
:
0
]
CAHBLTI0I1I
;
wire
[
31
:
0
]
CAHBLTl0I1I
;
wire
[
31
:
0
]
CAHBLTO1I1I
;
wire
[
31
:
0
]
CAHBLTI1I1I
;
wire
[
31
:
0
]
CAHBLTl1I1I
;
wire
[
31
:
0
]
CAHBLTOOl1I
;
wire
[
31
:
0
]
CAHBLTIOl1I
;
wire
[
31
:
0
]
CAHBLTlOl1I
;
wire
[
31
:
0
]
CAHBLTOIl1I
;
wire
[
31
:
0
]
CAHBLTO11l0
;
wire
[
31
:
0
]
CAHBLTI11l0
;
wire
[
31
:
0
]
CAHBLTl11l0
;
wire
[
31
:
0
]
CAHBLTOOO00
;
wire
[
31
:
0
]
CAHBLTIOO00
;
wire
[
31
:
0
]
CAHBLTlOO00
;
wire
[
31
:
0
]
CAHBLTOIO00
;
wire
[
31
:
0
]
CAHBLTIIO00
;
wire
[
31
:
0
]
CAHBLTlIO00
;
wire
[
31
:
0
]
CAHBLTOlO00
;
wire
[
31
:
0
]
CAHBLTIlO00
;
wire
[
31
:
0
]
CAHBLTllO00
;
wire
[
31
:
0
]
CAHBLTO0O00
;
wire
[
31
:
0
]
CAHBLTI0O00
;
wire
[
31
:
0
]
CAHBLTl0O00
;
wire
[
31
:
0
]
CAHBLTO1O00
;
wire
[
31
:
0
]
CAHBLTI1O00
;
wire
[
31
:
0
]
CAHBLTl1O00
;
wire
[
31
:
0
]
CAHBLTOOI00
;
wire
[
31
:
0
]
CAHBLTIOI00
;
wire
[
31
:
0
]
CAHBLTlOI00
;
wire
[
31
:
0
]
CAHBLTOII00
;
wire
[
31
:
0
]
CAHBLTIII00
;
wire
[
31
:
0
]
CAHBLTlII00
;
wire
[
31
:
0
]
CAHBLTOlI00
;
wire
[
31
:
0
]
CAHBLTIlI00
;
wire
[
31
:
0
]
CAHBLTllI00
;
wire
[
31
:
0
]
CAHBLTO0I00
;
wire
[
31
:
0
]
CAHBLTI0I00
;
wire
[
31
:
0
]
CAHBLTl0I00
;
wire
[
31
:
0
]
CAHBLTO1I00
;
wire
[
31
:
0
]
CAHBLTI1I00
;
wire
[
31
:
0
]
CAHBLTl1I00
;
wire
[
31
:
0
]
CAHBLTOOl00
;
wire
[
31
:
0
]
CAHBLTIIl1I
;
wire
[
31
:
0
]
CAHBLTlIl1I
;
wire
[
31
:
0
]
CAHBLTOll1I
;
wire
[
31
:
0
]
CAHBLTIll1I
;
wire
[
31
:
0
]
CAHBLTlll1I
;
wire
[
31
:
0
]
CAHBLTO0l1I
;
wire
[
31
:
0
]
CAHBLTI0l1I
;
wire
[
31
:
0
]
CAHBLTl0l1I
;
wire
[
31
:
0
]
CAHBLTO1l1I
;
wire
[
31
:
0
]
CAHBLTI1l1I
;
wire
[
31
:
0
]
CAHBLTl1l1I
;
wire
[
31
:
0
]
CAHBLTOO01I
;
wire
[
31
:
0
]
CAHBLTIO01I
;
wire
[
31
:
0
]
CAHBLTlO01I
;
wire
[
31
:
0
]
CAHBLTOI01I
;
wire
[
31
:
0
]
CAHBLTII01I
;
wire
[
31
:
0
]
CAHBLTlI01I
;
wire
[
31
:
0
]
CAHBLTOl01I
;
wire
[
31
:
0
]
CAHBLTIl01I
;
wire
[
31
:
0
]
CAHBLTll01I
;
wire
[
31
:
0
]
CAHBLTO001I
;
wire
[
31
:
0
]
CAHBLTI001I
;
wire
[
31
:
0
]
CAHBLTl001I
;
wire
[
31
:
0
]
CAHBLTO101I
;
wire
[
31
:
0
]
CAHBLTI101I
;
wire
[
31
:
0
]
CAHBLTl101I
;
wire
[
31
:
0
]
CAHBLTOO11I
;
wire
[
31
:
0
]
CAHBLTIO11I
;
wire
[
31
:
0
]
CAHBLTlO11I
;
wire
[
31
:
0
]
CAHBLTOI11I
;
wire
[
31
:
0
]
CAHBLTII11I
;
wire
[
31
:
0
]
CAHBLTlI11I
;
wire
[
31
:
0
]
CAHBLTOl11I
;
wire
[
31
:
0
]
CAHBLTIl11I
;
wire
[
31
:
0
]
CAHBLTIOl00
;
wire
[
31
:
0
]
CAHBLTlOl00
;
wire
[
31
:
0
]
CAHBLTOIl00
;
wire
[
31
:
0
]
CAHBLTIIl00
;
wire
[
31
:
0
]
CAHBLTlIl00
;
wire
[
31
:
0
]
CAHBLTOll00
;
wire
[
31
:
0
]
CAHBLTIll00
;
wire
[
31
:
0
]
CAHBLTlll00
;
wire
[
31
:
0
]
CAHBLTO0l00
;
wire
[
31
:
0
]
CAHBLTI0l00
;
wire
[
31
:
0
]
CAHBLTl0l00
;
wire
[
31
:
0
]
CAHBLTO1l00
;
wire
[
31
:
0
]
CAHBLTI1l00
;
wire
[
31
:
0
]
CAHBLTl1l00
;
wire
[
31
:
0
]
CAHBLTOO000
;
wire
[
31
:
0
]
CAHBLTIO000
;
wire
[
31
:
0
]
CAHBLTlO000
;
wire
[
31
:
0
]
CAHBLTOI000
;
wire
[
31
:
0
]
CAHBLTII000
;
wire
[
31
:
0
]
CAHBLTlI000
;
wire
[
31
:
0
]
CAHBLTOl000
;
wire
[
31
:
0
]
CAHBLTIl000
;
wire
[
31
:
0
]
CAHBLTll000
;
wire
[
31
:
0
]
CAHBLTO0000
;
wire
[
31
:
0
]
CAHBLTI0000
;
wire
[
31
:
0
]
CAHBLTl0000
;
wire
[
31
:
0
]
CAHBLTO1000
;
wire
[
31
:
0
]
CAHBLTI1000
;
wire
[
31
:
0
]
CAHBLTl1000
;
wire
[
31
:
0
]
CAHBLTOO100
;
wire
[
31
:
0
]
CAHBLTIO100
;
wire
[
31
:
0
]
CAHBLTlO100
;
wire
[
31
:
0
]
CAHBLTOI100
;
wire
[
31
:
0
]
CAHBLTII100
;
wire
[
2
:
0
]
CAHBLTll11I
;
wire
[
2
:
0
]
CAHBLTO011I
;
wire
[
2
:
0
]
CAHBLTI011I
;
wire
[
2
:
0
]
CAHBLTl011I
;
wire
[
2
:
0
]
CAHBLTO111I
;
wire
[
2
:
0
]
CAHBLTI111I
;
wire
[
2
:
0
]
CAHBLTl111I
;
wire
[
2
:
0
]
CAHBLTOOOOl
;
wire
[
2
:
0
]
CAHBLTIOOOl
;
wire
[
2
:
0
]
CAHBLTlOOOl
;
wire
[
2
:
0
]
CAHBLTOIOOl
;
wire
[
2
:
0
]
CAHBLTIIOOl
;
wire
[
2
:
0
]
CAHBLTlIOOl
;
wire
[
2
:
0
]
CAHBLTOlOOl
;
wire
[
2
:
0
]
CAHBLTIlOOl
;
wire
[
2
:
0
]
CAHBLTllOOl
;
wire
[
2
:
0
]
CAHBLTO0OOl
;
wire
[
2
:
0
]
CAHBLTI0OOl
;
wire
[
2
:
0
]
CAHBLTl0OOl
;
wire
[
2
:
0
]
CAHBLTO1OOl
;
wire
[
2
:
0
]
CAHBLTI1OOl
;
wire
[
2
:
0
]
CAHBLTl1OOl
;
wire
[
2
:
0
]
CAHBLTOOIOl
;
wire
[
2
:
0
]
CAHBLTIOIOl
;
wire
[
2
:
0
]
CAHBLTlOIOl
;
wire
[
2
:
0
]
CAHBLTOIIOl
;
wire
[
2
:
0
]
CAHBLTIIIOl
;
wire
[
2
:
0
]
CAHBLTlIIOl
;
wire
[
2
:
0
]
CAHBLTOlIOl
;
wire
[
2
:
0
]
CAHBLTIlIOl
;
wire
[
2
:
0
]
CAHBLTllIOl
;
wire
[
2
:
0
]
CAHBLTO0IOl
;
wire
[
2
:
0
]
CAHBLTI0IOl
;
wire
[
2
:
0
]
CAHBLTl0IOl
;
wire
[
2
:
0
]
CAHBLTlI100
;
wire
[
2
:
0
]
CAHBLTOl100
;
wire
[
2
:
0
]
CAHBLTIl100
;
wire
[
2
:
0
]
CAHBLTll100
;
wire
[
2
:
0
]
CAHBLTO0100
;
wire
[
2
:
0
]
CAHBLTI0100
;
wire
[
2
:
0
]
CAHBLTl0100
;
wire
[
2
:
0
]
CAHBLTO1100
;
wire
[
2
:
0
]
CAHBLTI1100
;
wire
[
2
:
0
]
CAHBLTl1100
;
wire
[
2
:
0
]
CAHBLTOOO10
;
wire
[
2
:
0
]
CAHBLTIOO10
;
wire
[
2
:
0
]
CAHBLTlOO10
;
wire
[
2
:
0
]
CAHBLTOIO10
;
wire
[
2
:
0
]
CAHBLTIIO10
;
wire
[
2
:
0
]
CAHBLTlIO10
;
wire
[
2
:
0
]
CAHBLTOlO10
;
wire
[
2
:
0
]
CAHBLTIlO10
;
wire
[
2
:
0
]
CAHBLTllO10
;
wire
[
2
:
0
]
CAHBLTO0O10
;
wire
[
2
:
0
]
CAHBLTI0O10
;
wire
[
2
:
0
]
CAHBLTl0O10
;
wire
[
2
:
0
]
CAHBLTO1O10
;
wire
[
2
:
0
]
CAHBLTI1O10
;
wire
[
2
:
0
]
CAHBLTl1O10
;
wire
[
2
:
0
]
CAHBLTOOI10
;
wire
[
2
:
0
]
CAHBLTIOI10
;
wire
[
2
:
0
]
CAHBLTlOI10
;
wire
[
2
:
0
]
CAHBLTOII10
;
wire
[
2
:
0
]
CAHBLTIII10
;
wire
[
2
:
0
]
CAHBLTlII10
;
wire
[
2
:
0
]
CAHBLTOlI10
;
wire
[
2
:
0
]
CAHBLTIlI10
;
wire
[
2
:
0
]
CAHBLTllI10
;
wire
CAHBLTO1IOl
;
wire
CAHBLTI1IOl
;
wire
CAHBLTl1IOl
;
wire
CAHBLTOOlOl
;
wire
CAHBLTIOlOl
;
wire
CAHBLTlOlOl
;
wire
CAHBLTOIlOl
;
wire
CAHBLTIIlOl
;
wire
CAHBLTlIlOl
;
wire
CAHBLTOllOl
;
wire
CAHBLTIllOl
;
wire
CAHBLTlllOl
;
wire
CAHBLTO0lOl
;
wire
CAHBLTI0lOl
;
wire
CAHBLTl0lOl
;
wire
CAHBLTO1lOl
;
wire
CAHBLTI1lOl
;
wire
CAHBLTl1lOl
;
wire
CAHBLTOO0Ol
;
wire
CAHBLTIO0Ol
;
wire
CAHBLTlO0Ol
;
wire
CAHBLTOI0Ol
;
wire
CAHBLTII0Ol
;
wire
CAHBLTlI0Ol
;
wire
CAHBLTOl0Ol
;
wire
CAHBLTIl0Ol
;
wire
CAHBLTll0Ol
;
wire
CAHBLTO00Ol
;
wire
CAHBLTI00Ol
;
wire
CAHBLTl00Ol
;
wire
CAHBLTO10Ol
;
wire
CAHBLTI10Ol
;
wire
CAHBLTl10Ol
;
wire
CAHBLTOO1Ol
;
wire
CAHBLTO0I10
;
wire
CAHBLTI0I10
;
wire
CAHBLTl0I10
;
wire
CAHBLTO1I10
;
wire
CAHBLTI1I10
;
wire
CAHBLTl1I10
;
wire
CAHBLTOOl10
;
wire
CAHBLTIOl10
;
wire
CAHBLTlOl10
;
wire
CAHBLTOIl10
;
wire
CAHBLTIIl10
;
wire
CAHBLTlIl10
;
wire
CAHBLTOll10
;
wire
CAHBLTIll10
;
wire
CAHBLTlll10
;
wire
CAHBLTO0l10
;
wire
CAHBLTI0l10
;
wire
CAHBLTl0l10
;
wire
CAHBLTO1l10
;
wire
CAHBLTI1l10
;
wire
CAHBLTl1l10
;
wire
CAHBLTOO010
;
wire
CAHBLTIO010
;
wire
CAHBLTlO010
;
wire
CAHBLTOI010
;
wire
CAHBLTII010
;
wire
CAHBLTlI010
;
wire
CAHBLTOl010
;
wire
CAHBLTIl010
;
wire
CAHBLTll010
;
wire
CAHBLTO0010
;
wire
CAHBLTI0010
;
wire
CAHBLTl0010
;
wire
CAHBLTO1010
;
wire
CAHBLTIO1Ol
;
wire
CAHBLTlO1Ol
;
wire
CAHBLTOI1Ol
;
wire
CAHBLTII1Ol
;
wire
CAHBLTlI1Ol
;
wire
CAHBLTOl1Ol
;
wire
CAHBLTIl1Ol
;
wire
CAHBLTll1Ol
;
wire
CAHBLTO01Ol
;
wire
CAHBLTI01Ol
;
wire
CAHBLTl01Ol
;
wire
CAHBLTO11Ol
;
wire
CAHBLTI11Ol
;
wire
CAHBLTl11Ol
;
wire
CAHBLTOOOIl
;
wire
CAHBLTIOOIl
;
wire
CAHBLTlOOIl
;
wire
CAHBLTOIOIl
;
wire
CAHBLTIIOIl
;
wire
CAHBLTlIOIl
;
wire
CAHBLTOlOIl
;
wire
CAHBLTIlOIl
;
wire
CAHBLTllOIl
;
wire
CAHBLTO0OIl
;
wire
CAHBLTI0OIl
;
wire
CAHBLTl0OIl
;
wire
CAHBLTO1OIl
;
wire
CAHBLTI1OIl
;
wire
CAHBLTl1OIl
;
wire
CAHBLTOOIIl
;
wire
CAHBLTIOIIl
;
wire
CAHBLTlOIIl
;
wire
CAHBLTOIIIl
;
wire
CAHBLTIIIIl
;
wire
CAHBLTI1010
;
wire
CAHBLTl1010
;
wire
CAHBLTOO110
;
wire
CAHBLTIO110
;
wire
CAHBLTlO110
;
wire
CAHBLTOI110
;
wire
CAHBLTII110
;
wire
CAHBLTlI110
;
wire
CAHBLTOl110
;
wire
CAHBLTIl110
;
wire
CAHBLTll110
;
wire
CAHBLTO0110
;
wire
CAHBLTI0110
;
wire
CAHBLTl0110
;
wire
CAHBLTO1110
;
wire
CAHBLTI1110
;
wire
CAHBLTl1110
;
wire
CAHBLTOOOO1
;
wire
CAHBLTIOOO1
;
wire
CAHBLTlOOO1
;
wire
CAHBLTOIOO1
;
wire
CAHBLTIIOO1
;
wire
CAHBLTlIOO1
;
wire
CAHBLTOlOO1
;
wire
CAHBLTIlOO1
;
wire
CAHBLTllOO1
;
wire
CAHBLTO0OO1
;
wire
CAHBLTI0OO1
;
wire
CAHBLTl0OO1
;
wire
CAHBLTO1OO1
;
wire
CAHBLTI1OO1
;
wire
CAHBLTl1OO1
;
wire
CAHBLTOOIO1
;
wire
CAHBLTIOIO1
;
wire
CAHBLTlIIIl
;
wire
CAHBLTOlIIl
;
wire
CAHBLTIlIIl
;
wire
CAHBLTllIIl
;
wire
CAHBLTO0IIl
;
wire
CAHBLTI0IIl
;
wire
CAHBLTl0IIl
;
wire
CAHBLTO1IIl
;
wire
CAHBLTI1IIl
;
wire
CAHBLTl1IIl
;
wire
CAHBLTOOlIl
;
wire
CAHBLTIOlIl
;
wire
CAHBLTlOlIl
;
wire
CAHBLTOIlIl
;
wire
CAHBLTIIlIl
;
wire
CAHBLTlIlIl
;
wire
CAHBLTOllIl
;
wire
CAHBLTIllIl
;
wire
CAHBLTlllIl
;
wire
CAHBLTO0lIl
;
wire
CAHBLTI0lIl
;
wire
CAHBLTl0lIl
;
wire
CAHBLTO1lIl
;
wire
CAHBLTI1lIl
;
wire
CAHBLTl1lIl
;
wire
CAHBLTOO0Il
;
wire
CAHBLTIO0Il
;
wire
CAHBLTlO0Il
;
wire
CAHBLTOI0Il
;
wire
CAHBLTII0Il
;
wire
CAHBLTlI0Il
;
wire
CAHBLTOl0Il
;
wire
CAHBLTIl0Il
;
wire
CAHBLTll0Il
;
wire
CAHBLTlOIO1
;
wire
CAHBLTOIIO1
;
wire
CAHBLTIIIO1
;
wire
CAHBLTlIIO1
;
wire
CAHBLTOlIO1
;
wire
CAHBLTIlIO1
;
wire
CAHBLTllIO1
;
wire
CAHBLTO0IO1
;
wire
CAHBLTI0IO1
;
wire
CAHBLTl0IO1
;
wire
CAHBLTO1IO1
;
wire
CAHBLTI1IO1
;
wire
CAHBLTl1IO1
;
wire
CAHBLTOOlO1
;
wire
CAHBLTIOlO1
;
wire
CAHBLTlOlO1
;
wire
CAHBLTOIlO1
;
wire
CAHBLTIIlO1
;
wire
CAHBLTlIlO1
;
wire
CAHBLTOllO1
;
wire
CAHBLTIllO1
;
wire
CAHBLTlllO1
;
wire
CAHBLTO0lO1
;
wire
CAHBLTI0lO1
;
wire
CAHBLTl0lO1
;
wire
CAHBLTO1lO1
;
wire
CAHBLTI1lO1
;
wire
CAHBLTl1lO1
;
wire
CAHBLTOO0O1
;
wire
CAHBLTIO0O1
;
wire
CAHBLTlO0O1
;
wire
CAHBLTOI0O1
;
wire
CAHBLTII0O1
;
wire
CAHBLTlI0O1
;
wire
CAHBLTO00Il
;
wire
CAHBLTI00Il
;
wire
CAHBLTl00Il
;
wire
CAHBLTO10Il
;
wire
CAHBLTI10Il
;
wire
CAHBLTl10Il
;
wire
CAHBLTOO1Il
;
wire
CAHBLTIO1Il
;
wire
CAHBLTlO1Il
;
wire
CAHBLTOI1Il
;
wire
CAHBLTII1Il
;
wire
CAHBLTlI1Il
;
wire
CAHBLTOl1Il
;
wire
CAHBLTIl1Il
;
wire
CAHBLTll1Il
;
wire
CAHBLTO01Il
;
wire
CAHBLTI01Il
;
wire
CAHBLTl01Il
;
wire
CAHBLTO11Il
;
wire
CAHBLTI11Il
;
wire
CAHBLTl11Il
;
wire
CAHBLTOOOll
;
wire
CAHBLTIOOll
;
wire
CAHBLTlOOll
;
wire
CAHBLTOIOll
;
wire
CAHBLTIIOll
;
wire
CAHBLTlIOll
;
wire
CAHBLTOlOll
;
wire
CAHBLTIlOll
;
wire
CAHBLTllOll
;
wire
CAHBLTO0Oll
;
wire
CAHBLTI0Oll
;
wire
CAHBLTl0Oll
;
wire
CAHBLTO1Oll
;
wire
CAHBLTOl0O1
;
wire
CAHBLTIl0O1
;
wire
CAHBLTll0O1
;
wire
CAHBLTO00O1
;
wire
CAHBLTI00O1
;
wire
CAHBLTl00O1
;
wire
CAHBLTO10O1
;
wire
CAHBLTI10O1
;
wire
CAHBLTl10O1
;
wire
CAHBLTOO1O1
;
wire
CAHBLTIO1O1
;
wire
CAHBLTlO1O1
;
wire
CAHBLTOI1O1
;
wire
CAHBLTII1O1
;
wire
CAHBLTlI1O1
;
wire
CAHBLTOl1O1
;
wire
CAHBLTIl1O1
;
wire
CAHBLTll1O1
;
wire
CAHBLTO01O1
;
wire
CAHBLTI01O1
;
wire
CAHBLTl01O1
;
wire
CAHBLTO11O1
;
wire
CAHBLTI11O1
;
wire
CAHBLTl11O1
;
wire
CAHBLTOOOI1
;
wire
CAHBLTIOOI1
;
wire
CAHBLTlOOI1
;
wire
CAHBLTOIOI1
;
wire
CAHBLTIIOI1
;
wire
CAHBLTlIOI1
;
wire
CAHBLTOlOI1
;
wire
CAHBLTIlOI1
;
wire
CAHBLTllOI1
;
wire
CAHBLTO0OI1
;
wire
CAHBLTI1Oll
;
wire
CAHBLTl1Oll
;
wire
CAHBLTI0OI1
;
wire
CAHBLTl0OI1
;
generate
if
(
CAHBLTIIO0
[
0
]
)
assign
CAHBLTl1O0
=
CAHBLTO0O0
;
else
assign
CAHBLTl1O0
=
1
'b
1
;
if
(
CAHBLTIIO0
[
1
]
)
assign
CAHBLTO0I0
=
CAHBLTIII0
;
else
assign
CAHBLTO0I0
=
1
'b
1
;
if
(
CAHBLTIIO0
[
2
]
)
assign
CAHBLTIIl0
=
CAHBLTl1I0
;
else
assign
CAHBLTIIl0
=
1
'b
1
;
if
(
CAHBLTIIO0
[
3
]
)
assign
CAHBLTl1l0
=
CAHBLTO0l0
;
else
assign
CAHBLTl1l0
=
1
'b
1
;
if
(
CAHBLTIIO0
[
4
]
)
assign
CAHBLTO000
=
CAHBLTII00
;
else
assign
CAHBLTO000
=
1
'b
1
;
if
(
CAHBLTIIO0
[
5
]
)
assign
CAHBLTII10
=
CAHBLTl100
;
else
assign
CAHBLTII10
=
1
'b
1
;
if
(
CAHBLTIIO0
[
6
]
)
assign
CAHBLTl110
=
CAHBLTO010
;
else
assign
CAHBLTl110
=
1
'b
1
;
if
(
CAHBLTIIO0
[
7
]
)
assign
CAHBLTO0O1
=
CAHBLTIIO1
;
else
assign
CAHBLTO0O1
=
1
'b
1
;
if
(
CAHBLTIIO0
[
8
]
)
assign
CAHBLTIII1
=
CAHBLTl1O1
;
else
assign
CAHBLTIII1
=
1
'b
1
;
if
(
CAHBLTIIO0
[
9
]
)
assign
CAHBLTl1I1
=
CAHBLTO0I1
;
else
assign
CAHBLTl1I1
=
1
'b
1
;
if
(
CAHBLTIIO0
[
10
]
)
assign
CAHBLTO0l1
=
CAHBLTIIl1
;
else
assign
CAHBLTO0l1
=
1
'b
1
;
if
(
CAHBLTIIO0
[
11
]
)
assign
CAHBLTII01
=
CAHBLTl1l1
;
else
assign
CAHBLTII01
=
1
'b
1
;
if
(
CAHBLTIIO0
[
12
]
)
assign
CAHBLTl101
=
CAHBLTO001
;
else
assign
CAHBLTl101
=
1
'b
1
;
if
(
CAHBLTIIO0
[
13
]
)
assign
CAHBLTO011
=
CAHBLTII11
;
else
assign
CAHBLTO011
=
1
'b
1
;
if
(
CAHBLTIIO0
[
14
]
)
assign
CAHBLTIIOOI
=
CAHBLTl111
;
else
assign
CAHBLTIIOOI
=
1
'b
1
;
if
(
CAHBLTIIO0
[
15
]
)
assign
CAHBLTl1OOI
=
CAHBLTO0OOI
;
else
assign
CAHBLTl1OOI
=
1
'b
1
;
if
(
CAHBLTIIO0
[
16
]
)
assign
CAHBLTO0IOI
=
CAHBLTIIIOI
;
else
assign
CAHBLTO0IOI
=
1
'b
1
;
if
(
CAHBLTlIO0
[
0
]
)
assign
CAHBLTlIlOI
=
CAHBLTOOlOI
;
else
assign
CAHBLTlIlOI
=
1
'b
1
;
if
(
CAHBLTlIO0
[
1
]
)
assign
CAHBLTOO0OI
=
CAHBLTI0lOI
;
else
assign
CAHBLTOO0OI
=
1
'b
1
;
if
(
CAHBLTlIO0
[
2
]
)
assign
CAHBLTI00OI
=
CAHBLTlI0OI
;
else
assign
CAHBLTI00OI
=
1
'b
1
;
if
(
CAHBLTlIO0
[
3
]
)
assign
CAHBLTlI1OI
=
CAHBLTOO1OI
;
else
assign
CAHBLTlI1OI
=
1
'b
1
;
if
(
CAHBLTlIO0
[
4
]
)
assign
CAHBLTOOOII
=
CAHBLTI01OI
;
else
assign
CAHBLTOOOII
=
1
'b
1
;
if
(
CAHBLTlIO0
[
5
]
)
assign
CAHBLTI0OII
=
CAHBLTlIOII
;
else
assign
CAHBLTI0OII
=
1
'b
1
;
if
(
CAHBLTlIO0
[
6
]
)
assign
CAHBLTlIIII
=
CAHBLTOOIII
;
else
assign
CAHBLTlIIII
=
1
'b
1
;
if
(
CAHBLTlIO0
[
7
]
)
assign
CAHBLTOOlII
=
CAHBLTI0III
;
else
assign
CAHBLTOOlII
=
1
'b
1
;
if
(
CAHBLTlIO0
[
8
]
)
assign
CAHBLTI0lII
=
CAHBLTlIlII
;
else
assign
CAHBLTI0lII
=
1
'b
1
;
if
(
CAHBLTlIO0
[
9
]
)
assign
CAHBLTlI0II
=
CAHBLTOO0II
;
else
assign
CAHBLTlI0II
=
1
'b
1
;
if
(
CAHBLTlIO0
[
10
]
)
assign
CAHBLTOO1II
=
CAHBLTI00II
;
else
assign
CAHBLTOO1II
=
1
'b
1
;
if
(
CAHBLTlIO0
[
11
]
)
assign
CAHBLTI01II
=
CAHBLTlI1II
;
else
assign
CAHBLTI01II
=
1
'b
1
;
if
(
CAHBLTlIO0
[
12
]
)
assign
CAHBLTlIOlI
=
CAHBLTOOOlI
;
else
assign
CAHBLTlIOlI
=
1
'b
1
;
if
(
CAHBLTlIO0
[
13
]
)
assign
CAHBLTOOIlI
=
CAHBLTI0OlI
;
else
assign
CAHBLTOOIlI
=
1
'b
1
;
if
(
CAHBLTlIO0
[
14
]
)
assign
CAHBLTI0IlI
=
CAHBLTlIIlI
;
else
assign
CAHBLTI0IlI
=
1
'b
1
;
if
(
CAHBLTlIO0
[
15
]
)
assign
CAHBLTlIllI
=
CAHBLTOOllI
;
else
assign
CAHBLTlIllI
=
1
'b
1
;
if
(
CAHBLTlIO0
[
16
]
)
assign
CAHBLTOO0lI
=
CAHBLTI0llI
;
else
assign
CAHBLTOO0lI
=
1
'b
1
;
if
(
CAHBLTlIlll
[
0
]
)
assign
CAHBLTOO0ll
=
CAHBLTI0lll
;
else
assign
CAHBLTOO0ll
=
1
'b
1
;
if
(
CAHBLTlIlll
[
1
]
)
assign
CAHBLTI00ll
=
CAHBLTlI0ll
;
else
assign
CAHBLTI00ll
=
1
'b
1
;
if
(
CAHBLTlIlll
[
2
]
)
assign
CAHBLTlI1ll
=
CAHBLTOO1ll
;
else
assign
CAHBLTlI1ll
=
1
'b
1
;
if
(
CAHBLTlIlll
[
3
]
)
assign
CAHBLTOOO0l
=
CAHBLTI01ll
;
else
assign
CAHBLTOOO0l
=
1
'b
1
;
if
(
CAHBLTlIlll
[
4
]
)
assign
CAHBLTI0O0l
=
CAHBLTlIO0l
;
else
assign
CAHBLTI0O0l
=
1
'b
1
;
if
(
CAHBLTlIlll
[
5
]
)
assign
CAHBLTlII0l
=
CAHBLTOOI0l
;
else
assign
CAHBLTlII0l
=
1
'b
1
;
if
(
CAHBLTlIlll
[
6
]
)
assign
CAHBLTOOl0l
=
CAHBLTI0I0l
;
else
assign
CAHBLTOOl0l
=
1
'b
1
;
if
(
CAHBLTlIlll
[
7
]
)
assign
CAHBLTI0l0l
=
CAHBLTlIl0l
;
else
assign
CAHBLTI0l0l
=
1
'b
1
;
if
(
CAHBLTlIlll
[
8
]
)
assign
CAHBLTlI00l
=
CAHBLTOO00l
;
else
assign
CAHBLTlI00l
=
1
'b
1
;
if
(
CAHBLTlIlll
[
9
]
)
assign
CAHBLTOO10l
=
CAHBLTI000l
;
else
assign
CAHBLTOO10l
=
1
'b
1
;
if
(
CAHBLTlIlll
[
10
]
)
assign
CAHBLTI010l
=
CAHBLTlI10l
;
else
assign
CAHBLTI010l
=
1
'b
1
;
if
(
CAHBLTlIlll
[
11
]
)
assign
CAHBLTlIO1l
=
CAHBLTOOO1l
;
else
assign
CAHBLTlIO1l
=
1
'b
1
;
if
(
CAHBLTlIlll
[
12
]
)
assign
CAHBLTOOI1l
=
CAHBLTI0O1l
;
else
assign
CAHBLTOOI1l
=
1
'b
1
;
if
(
CAHBLTlIlll
[
13
]
)
assign
CAHBLTI0I1l
=
CAHBLTlII1l
;
else
assign
CAHBLTI0I1l
=
1
'b
1
;
if
(
CAHBLTlIlll
[
14
]
)
assign
CAHBLTlIl1l
=
CAHBLTOOl1l
;
else
assign
CAHBLTlIl1l
=
1
'b
1
;
if
(
CAHBLTlIlll
[
15
]
)
assign
CAHBLTOO01l
=
CAHBLTI0l1l
;
else
assign
CAHBLTOO01l
=
1
'b
1
;
if
(
CAHBLTlIlll
[
16
]
)
assign
CAHBLTI001l
=
CAHBLTlI01l
;
else
assign
CAHBLTI001l
=
1
'b
1
;
if
(
CAHBLTOllll
[
0
]
)
assign
CAHBLTOl11l
=
CAHBLTIO11l
;
else
assign
CAHBLTOl11l
=
1
'b
1
;
if
(
CAHBLTOllll
[
1
]
)
assign
CAHBLTIOOO0
=
CAHBLTl011l
;
else
assign
CAHBLTIOOO0
=
1
'b
1
;
if
(
CAHBLTOllll
[
2
]
)
assign
CAHBLTl0OO0
=
CAHBLTOlOO0
;
else
assign
CAHBLTl0OO0
=
1
'b
1
;
if
(
CAHBLTOllll
[
3
]
)
assign
CAHBLTOlIO0
=
CAHBLTIOIO0
;
else
assign
CAHBLTOlIO0
=
1
'b
1
;
if
(
CAHBLTOllll
[
4
]
)
assign
CAHBLTIOlO0
=
CAHBLTl0IO0
;
else
assign
CAHBLTIOlO0
=
1
'b
1
;
if
(
CAHBLTOllll
[
5
]
)
assign
CAHBLTl0lO0
=
CAHBLTOllO0
;
else
assign
CAHBLTl0lO0
=
1
'b
1
;
if
(
CAHBLTOllll
[
6
]
)
assign
CAHBLTOl0O0
=
CAHBLTIO0O0
;
else
assign
CAHBLTOl0O0
=
1
'b
1
;
if
(
CAHBLTOllll
[
7
]
)
assign
CAHBLTIO1O0
=
CAHBLTl00O0
;
else
assign
CAHBLTIO1O0
=
1
'b
1
;
if
(
CAHBLTOllll
[
8
]
)
assign
CAHBLTl01O0
=
CAHBLTOl1O0
;
else
assign
CAHBLTl01O0
=
1
'b
1
;
if
(
CAHBLTOllll
[
9
]
)
assign
CAHBLTOlOI0
=
CAHBLTIOOI0
;
else
assign
CAHBLTOlOI0
=
1
'b
1
;
if
(
CAHBLTOllll
[
10
]
)
assign
CAHBLTIOII0
=
CAHBLTl0OI0
;
else
assign
CAHBLTIOII0
=
1
'b
1
;
if
(
CAHBLTOllll
[
11
]
)
assign
CAHBLTl0II0
=
CAHBLTOlII0
;
else
assign
CAHBLTl0II0
=
1
'b
1
;
if
(
CAHBLTOllll
[
12
]
)
assign
CAHBLTOllI0
=
CAHBLTIOlI0
;
else
assign
CAHBLTOllI0
=
1
'b
1
;
if
(
CAHBLTOllll
[
13
]
)
assign
CAHBLTIO0I0
=
CAHBLTl0lI0
;
else
assign
CAHBLTIO0I0
=
1
'b
1
;
if
(
CAHBLTOllll
[
14
]
)
assign
CAHBLTl00I0
=
CAHBLTOl0I0
;
else
assign
CAHBLTl00I0
=
1
'b
1
;
if
(
CAHBLTOllll
[
15
]
)
assign
CAHBLTOl1I0
=
CAHBLTIO1I0
;
else
assign
CAHBLTOl1I0
=
1
'b
1
;
if
(
CAHBLTOllll
[
16
]
)
assign
CAHBLTIOOl0
=
CAHBLTl01I0
;
else
assign
CAHBLTIOOl0
=
1
'b
1
;
endgenerate
generate
if
(
CAHBLTIIO0
[
0
]
)
assign
CAHBLTOOI0
=
CAHBLTI0O0
;
else
assign
CAHBLTOOI0
=
1
'b
1
;
if
(
CAHBLTIIO0
[
1
]
)
assign
CAHBLTI0I0
=
CAHBLTlII0
;
else
assign
CAHBLTI0I0
=
1
'b
1
;
if
(
CAHBLTIIO0
[
2
]
)
assign
CAHBLTlIl0
=
CAHBLTOOl0
;
else
assign
CAHBLTlIl0
=
1
'b
1
;
if
(
CAHBLTIIO0
[
3
]
)
assign
CAHBLTOO00
=
CAHBLTI0l0
;
else
assign
CAHBLTOO00
=
1
'b
1
;
if
(
CAHBLTIIO0
[
4
]
)
assign
CAHBLTI000
=
CAHBLTlI00
;
else
assign
CAHBLTI000
=
1
'b
1
;
if
(
CAHBLTIIO0
[
5
]
)
assign
CAHBLTlI10
=
CAHBLTOO10
;
else
assign
CAHBLTlI10
=
1
'b
1
;
if
(
CAHBLTIIO0
[
6
]
)
assign
CAHBLTOOO1
=
CAHBLTI010
;
else
assign
CAHBLTOOO1
=
1
'b
1
;
if
(
CAHBLTIIO0
[
7
]
)
assign
CAHBLTI0O1
=
CAHBLTlIO1
;
else
assign
CAHBLTI0O1
=
1
'b
1
;
if
(
CAHBLTIIO0
[
8
]
)
assign
CAHBLTlII1
=
CAHBLTOOI1
;
else
assign
CAHBLTlII1
=
1
'b
1
;
if
(
CAHBLTIIO0
[
9
]
)
assign
CAHBLTOOl1
=
CAHBLTI0I1
;
else
assign
CAHBLTOOl1
=
1
'b
1
;
if
(
CAHBLTIIO0
[
10
]
)
assign
CAHBLTI0l1
=
CAHBLTlIl1
;
else
assign
CAHBLTI0l1
=
1
'b
1
;
if
(
CAHBLTIIO0
[
11
]
)
assign
CAHBLTlI01
=
CAHBLTOO01
;
else
assign
CAHBLTlI01
=
1
'b
1
;
if
(
CAHBLTIIO0
[
12
]
)
assign
CAHBLTOO11
=
CAHBLTI001
;
else
assign
CAHBLTOO11
=
1
'b
1
;
if
(
CAHBLTIIO0
[
13
]
)
assign
CAHBLTI011
=
CAHBLTlI11
;
else
assign
CAHBLTI011
=
1
'b
1
;
if
(
CAHBLTIIO0
[
14
]
)
assign
CAHBLTlIOOI
=
CAHBLTOOOOI
;
else
assign
CAHBLTlIOOI
=
1
'b
1
;
if
(
CAHBLTIIO0
[
15
]
)
assign
CAHBLTOOIOI
=
CAHBLTI0OOI
;
else
assign
CAHBLTOOIOI
=
1
'b
1
;
if
(
CAHBLTIIO0
[
16
]
)
assign
CAHBLTI0IOI
=
CAHBLTlIIOI
;
else
assign
CAHBLTI0IOI
=
1
'b
1
;
if
(
CAHBLTlIO0
[
0
]
)
assign
CAHBLTOllOI
=
CAHBLTIOlOI
;
else
assign
CAHBLTOllOI
=
1
'b
1
;
if
(
CAHBLTlIO0
[
1
]
)
assign
CAHBLTIO0OI
=
CAHBLTl0lOI
;
else
assign
CAHBLTIO0OI
=
1
'b
1
;
if
(
CAHBLTlIO0
[
2
]
)
assign
CAHBLTl00OI
=
CAHBLTOl0OI
;
else
assign
CAHBLTl00OI
=
1
'b
1
;
if
(
CAHBLTlIO0
[
3
]
)
assign
CAHBLTOl1OI
=
CAHBLTIO1OI
;
else
assign
CAHBLTOl1OI
=
1
'b
1
;
if
(
CAHBLTlIO0
[
4
]
)
assign
CAHBLTIOOII
=
CAHBLTl01OI
;
else
assign
CAHBLTIOOII
=
1
'b
1
;
if
(
CAHBLTlIO0
[
5
]
)
assign
CAHBLTl0OII
=
CAHBLTOlOII
;
else
assign
CAHBLTl0OII
=
1
'b
1
;
if
(
CAHBLTlIO0
[
6
]
)
assign
CAHBLTOlIII
=
CAHBLTIOIII
;
else
assign
CAHBLTOlIII
=
1
'b
1
;
if
(
CAHBLTlIO0
[
7
]
)
assign
CAHBLTIOlII
=
CAHBLTl0III
;
else
assign
CAHBLTIOlII
=
1
'b
1
;
if
(
CAHBLTlIO0
[
8
]
)
assign
CAHBLTl0lII
=
CAHBLTOllII
;
else
assign
CAHBLTl0lII
=
1
'b
1
;
if
(
CAHBLTlIO0
[
9
]
)
assign
CAHBLTOl0II
=
CAHBLTIO0II
;
else
assign
CAHBLTOl0II
=
1
'b
1
;
if
(
CAHBLTlIO0
[
10
]
)
assign
CAHBLTIO1II
=
CAHBLTl00II
;
else
assign
CAHBLTIO1II
=
1
'b
1
;
if
(
CAHBLTlIO0
[
11
]
)
assign
CAHBLTl01II
=
CAHBLTOl1II
;
else
assign
CAHBLTl01II
=
1
'b
1
;
if
(
CAHBLTlIO0
[
12
]
)
assign
CAHBLTOlOlI
=
CAHBLTIOOlI
;
else
assign
CAHBLTOlOlI
=
1
'b
1
;
if
(
CAHBLTlIO0
[
13
]
)
assign
CAHBLTIOIlI
=
CAHBLTl0OlI
;
else
assign
CAHBLTIOIlI
=
1
'b
1
;
if
(
CAHBLTlIO0
[
14
]
)
assign
CAHBLTl0IlI
=
CAHBLTOlIlI
;
else
assign
CAHBLTl0IlI
=
1
'b
1
;
if
(
CAHBLTlIO0
[
15
]
)
assign
CAHBLTOlllI
=
CAHBLTIOllI
;
else
assign
CAHBLTOlllI
=
1
'b
1
;
if
(
CAHBLTlIO0
[
16
]
)
assign
CAHBLTIO0lI
=
CAHBLTl0llI
;
else
assign
CAHBLTIO0lI
=
1
'b
1
;
if
(
CAHBLTlIlll
[
0
]
)
assign
CAHBLTIO0ll
=
CAHBLTl0lll
;
else
assign
CAHBLTIO0ll
=
1
'b
1
;
if
(
CAHBLTlIlll
[
1
]
)
assign
CAHBLTl00ll
=
CAHBLTOl0ll
;
else
assign
CAHBLTl00ll
=
1
'b
1
;
if
(
CAHBLTlIlll
[
2
]
)
assign
CAHBLTOl1ll
=
CAHBLTIO1ll
;
else
assign
CAHBLTOl1ll
=
1
'b
1
;
if
(
CAHBLTlIlll
[
3
]
)
assign
CAHBLTIOO0l
=
CAHBLTl01ll
;
else
assign
CAHBLTIOO0l
=
1
'b
1
;
if
(
CAHBLTlIlll
[
4
]
)
assign
CAHBLTl0O0l
=
CAHBLTOlO0l
;
else
assign
CAHBLTl0O0l
=
1
'b
1
;
if
(
CAHBLTlIlll
[
5
]
)
assign
CAHBLTOlI0l
=
CAHBLTIOI0l
;
else
assign
CAHBLTOlI0l
=
1
'b
1
;
if
(
CAHBLTlIlll
[
6
]
)
assign
CAHBLTIOl0l
=
CAHBLTl0I0l
;
else
assign
CAHBLTIOl0l
=
1
'b
1
;
if
(
CAHBLTlIlll
[
7
]
)
assign
CAHBLTl0l0l
=
CAHBLTOll0l
;
else
assign
CAHBLTl0l0l
=
1
'b
1
;
if
(
CAHBLTlIlll
[
8
]
)
assign
CAHBLTOl00l
=
CAHBLTIO00l
;
else
assign
CAHBLTOl00l
=
1
'b
1
;
if
(
CAHBLTlIlll
[
9
]
)
assign
CAHBLTIO10l
=
CAHBLTl000l
;
else
assign
CAHBLTIO10l
=
1
'b
1
;
if
(
CAHBLTlIlll
[
10
]
)
assign
CAHBLTl010l
=
CAHBLTOl10l
;
else
assign
CAHBLTl010l
=
1
'b
1
;
if
(
CAHBLTlIlll
[
11
]
)
assign
CAHBLTOlO1l
=
CAHBLTIOO1l
;
else
assign
CAHBLTOlO1l
=
1
'b
1
;
if
(
CAHBLTlIlll
[
12
]
)
assign
CAHBLTIOI1l
=
CAHBLTl0O1l
;
else
assign
CAHBLTIOI1l
=
1
'b
1
;
if
(
CAHBLTlIlll
[
13
]
)
assign
CAHBLTl0I1l
=
CAHBLTOlI1l
;
else
assign
CAHBLTl0I1l
=
1
'b
1
;
if
(
CAHBLTlIlll
[
14
]
)
assign
CAHBLTOll1l
=
CAHBLTIOl1l
;
else
assign
CAHBLTOll1l
=
1
'b
1
;
if
(
CAHBLTlIlll
[
15
]
)
assign
CAHBLTIO01l
=
CAHBLTl0l1l
;
else
assign
CAHBLTIO01l
=
1
'b
1
;
if
(
CAHBLTlIlll
[
16
]
)
assign
CAHBLTl001l
=
CAHBLTOl01l
;
else
assign
CAHBLTl001l
=
1
'b
1
;
if
(
CAHBLTOllll
[
0
]
)
assign
CAHBLTIl11l
=
CAHBLTlO11l
;
else
assign
CAHBLTIl11l
=
1
'b
1
;
if
(
CAHBLTOllll
[
1
]
)
assign
CAHBLTlOOO0
=
CAHBLTO111l
;
else
assign
CAHBLTlOOO0
=
1
'b
1
;
if
(
CAHBLTOllll
[
2
]
)
assign
CAHBLTO1OO0
=
CAHBLTIlOO0
;
else
assign
CAHBLTO1OO0
=
1
'b
1
;
if
(
CAHBLTOllll
[
3
]
)
assign
CAHBLTIlIO0
=
CAHBLTlOIO0
;
else
assign
CAHBLTIlIO0
=
1
'b
1
;
if
(
CAHBLTOllll
[
4
]
)
assign
CAHBLTlOlO0
=
CAHBLTO1IO0
;
else
assign
CAHBLTlOlO0
=
1
'b
1
;
if
(
CAHBLTOllll
[
5
]
)
assign
CAHBLTO1lO0
=
CAHBLTIllO0
;
else
assign
CAHBLTO1lO0
=
1
'b
1
;
if
(
CAHBLTOllll
[
6
]
)
assign
CAHBLTIl0O0
=
CAHBLTlO0O0
;
else
assign
CAHBLTIl0O0
=
1
'b
1
;
if
(
CAHBLTOllll
[
7
]
)
assign
CAHBLTlO1O0
=
CAHBLTO10O0
;
else
assign
CAHBLTlO1O0
=
1
'b
1
;
if
(
CAHBLTOllll
[
8
]
)
assign
CAHBLTO11O0
=
CAHBLTIl1O0
;
else
assign
CAHBLTO11O0
=
1
'b
1
;
if
(
CAHBLTOllll
[
9
]
)
assign
CAHBLTIlOI0
=
CAHBLTlOOI0
;
else
assign
CAHBLTIlOI0
=
1
'b
1
;
if
(
CAHBLTOllll
[
10
]
)
assign
CAHBLTlOII0
=
CAHBLTO1OI0
;
else
assign
CAHBLTlOII0
=
1
'b
1
;
if
(
CAHBLTOllll
[
11
]
)
assign
CAHBLTO1II0
=
CAHBLTIlII0
;
else
assign
CAHBLTO1II0
=
1
'b
1
;
if
(
CAHBLTOllll
[
12
]
)
assign
CAHBLTIllI0
=
CAHBLTlOlI0
;
else
assign
CAHBLTIllI0
=
1
'b
1
;
if
(
CAHBLTOllll
[
13
]
)
assign
CAHBLTlO0I0
=
CAHBLTO1lI0
;
else
assign
CAHBLTlO0I0
=
1
'b
1
;
if
(
CAHBLTOllll
[
14
]
)
assign
CAHBLTO10I0
=
CAHBLTIl0I0
;
else
assign
CAHBLTO10I0
=
1
'b
1
;
if
(
CAHBLTOllll
[
15
]
)
assign
CAHBLTIl1I0
=
CAHBLTlO1I0
;
else
assign
CAHBLTIl1I0
=
1
'b
1
;
if
(
CAHBLTOllll
[
16
]
)
assign
CAHBLTlOOl0
=
CAHBLTO11I0
;
else
assign
CAHBLTlOOl0
=
1
'b
1
;
endgenerate
generate
if
(
CAHBLTIIO0
[
0
]
)
assign
CAHBLTIOI0
=
CAHBLTl0O0
;
else
assign
CAHBLTIOI0
=
1
'b
0
;
if
(
CAHBLTIIO0
[
1
]
)
assign
CAHBLTl0I0
=
CAHBLTOlI0
;
else
assign
CAHBLTl0I0
=
1
'b
0
;
if
(
CAHBLTIIO0
[
2
]
)
assign
CAHBLTOll0
=
CAHBLTIOl0
;
else
assign
CAHBLTOll0
=
1
'b
0
;
if
(
CAHBLTIIO0
[
3
]
)
assign
CAHBLTIO00
=
CAHBLTl0l0
;
else
assign
CAHBLTIO00
=
1
'b
0
;
if
(
CAHBLTIIO0
[
4
]
)
assign
CAHBLTl000
=
CAHBLTOl00
;
else
assign
CAHBLTl000
=
1
'b
0
;
if
(
CAHBLTIIO0
[
5
]
)
assign
CAHBLTOl10
=
CAHBLTIO10
;
else
assign
CAHBLTOl10
=
1
'b
0
;
if
(
CAHBLTIIO0
[
6
]
)
assign
CAHBLTIOO1
=
CAHBLTl010
;
else
assign
CAHBLTIOO1
=
1
'b
0
;
if
(
CAHBLTIIO0
[
7
]
)
assign
CAHBLTl0O1
=
CAHBLTOlO1
;
else
assign
CAHBLTl0O1
=
1
'b
0
;
if
(
CAHBLTIIO0
[
8
]
)
assign
CAHBLTOlI1
=
CAHBLTIOI1
;
else
assign
CAHBLTOlI1
=
1
'b
0
;
if
(
CAHBLTIIO0
[
9
]
)
assign
CAHBLTIOl1
=
CAHBLTl0I1
;
else
assign
CAHBLTIOl1
=
1
'b
0
;
if
(
CAHBLTIIO0
[
10
]
)
assign
CAHBLTl0l1
=
CAHBLTOll1
;
else
assign
CAHBLTl0l1
=
1
'b
0
;
if
(
CAHBLTIIO0
[
11
]
)
assign
CAHBLTOl01
=
CAHBLTIO01
;
else
assign
CAHBLTOl01
=
1
'b
0
;
if
(
CAHBLTIIO0
[
12
]
)
assign
CAHBLTIO11
=
CAHBLTl001
;
else
assign
CAHBLTIO11
=
1
'b
0
;
if
(
CAHBLTIIO0
[
13
]
)
assign
CAHBLTl011
=
CAHBLTOl11
;
else
assign
CAHBLTl011
=
1
'b
0
;
if
(
CAHBLTIIO0
[
14
]
)
assign
CAHBLTOlOOI
=
CAHBLTIOOOI
;
else
assign
CAHBLTOlOOI
=
1
'b
0
;
if
(
CAHBLTIIO0
[
15
]
)
assign
CAHBLTIOIOI
=
CAHBLTl0OOI
;
else
assign
CAHBLTIOIOI
=
1
'b
0
;
if
(
CAHBLTIIO0
[
16
]
)
assign
CAHBLTl0IOI
=
CAHBLTOlIOI
;
else
assign
CAHBLTl0IOI
=
1
'b
0
;
if
(
CAHBLTlIO0
[
0
]
)
assign
CAHBLTIllOI
=
CAHBLTlOlOI
;
else
assign
CAHBLTIllOI
=
1
'b
0
;
if
(
CAHBLTlIO0
[
1
]
)
assign
CAHBLTlO0OI
=
CAHBLTO1lOI
;
else
assign
CAHBLTlO0OI
=
1
'b
0
;
if
(
CAHBLTlIO0
[
2
]
)
assign
CAHBLTO10OI
=
CAHBLTIl0OI
;
else
assign
CAHBLTO10OI
=
1
'b
0
;
if
(
CAHBLTlIO0
[
3
]
)
assign
CAHBLTIl1OI
=
CAHBLTlO1OI
;
else
assign
CAHBLTIl1OI
=
1
'b
0
;
if
(
CAHBLTlIO0
[
4
]
)
assign
CAHBLTlOOII
=
CAHBLTO11OI
;
else
assign
CAHBLTlOOII
=
1
'b
0
;
if
(
CAHBLTlIO0
[
5
]
)
assign
CAHBLTO1OII
=
CAHBLTIlOII
;
else
assign
CAHBLTO1OII
=
1
'b
0
;
if
(
CAHBLTlIO0
[
6
]
)
assign
CAHBLTIlIII
=
CAHBLTlOIII
;
else
assign
CAHBLTIlIII
=
1
'b
0
;
if
(
CAHBLTlIO0
[
7
]
)
assign
CAHBLTlOlII
=
CAHBLTO1III
;
else
assign
CAHBLTlOlII
=
1
'b
0
;
if
(
CAHBLTlIO0
[
8
]
)
assign
CAHBLTO1lII
=
CAHBLTIllII
;
else
assign
CAHBLTO1lII
=
1
'b
0
;
if
(
CAHBLTlIO0
[
9
]
)
assign
CAHBLTIl0II
=
CAHBLTlO0II
;
else
assign
CAHBLTIl0II
=
1
'b
0
;
if
(
CAHBLTlIO0
[
10
]
)
assign
CAHBLTlO1II
=
CAHBLTO10II
;
else
assign
CAHBLTlO1II
=
1
'b
0
;
if
(
CAHBLTlIO0
[
11
]
)
assign
CAHBLTO11II
=
CAHBLTIl1II
;
else
assign
CAHBLTO11II
=
1
'b
0
;
if
(
CAHBLTlIO0
[
12
]
)
assign
CAHBLTIlOlI
=
CAHBLTlOOlI
;
else
assign
CAHBLTIlOlI
=
1
'b
0
;
if
(
CAHBLTlIO0
[
13
]
)
assign
CAHBLTlOIlI
=
CAHBLTO1OlI
;
else
assign
CAHBLTlOIlI
=
1
'b
0
;
if
(
CAHBLTlIO0
[
14
]
)
assign
CAHBLTO1IlI
=
CAHBLTIlIlI
;
else
assign
CAHBLTO1IlI
=
1
'b
0
;
if
(
CAHBLTlIO0
[
15
]
)
assign
CAHBLTIlllI
=
CAHBLTlOllI
;
else
assign
CAHBLTIlllI
=
1
'b
0
;
if
(
CAHBLTlIO0
[
16
]
)
assign
CAHBLTlO0lI
=
CAHBLTO1llI
;
else
assign
CAHBLTlO0lI
=
1
'b
0
;
if
(
CAHBLTlIlll
[
0
]
)
assign
CAHBLTlO0ll
=
CAHBLTO1lll
;
else
assign
CAHBLTlO0ll
=
1
'b
0
;
if
(
CAHBLTlIlll
[
1
]
)
assign
CAHBLTO10ll
=
CAHBLTIl0ll
;
else
assign
CAHBLTO10ll
=
1
'b
0
;
if
(
CAHBLTlIlll
[
2
]
)
assign
CAHBLTIl1ll
=
CAHBLTlO1ll
;
else
assign
CAHBLTIl1ll
=
1
'b
0
;
if
(
CAHBLTlIlll
[
3
]
)
assign
CAHBLTlOO0l
=
CAHBLTO11ll
;
else
assign
CAHBLTlOO0l
=
1
'b
0
;
if
(
CAHBLTlIlll
[
4
]
)
assign
CAHBLTO1O0l
=
CAHBLTIlO0l
;
else
assign
CAHBLTO1O0l
=
1
'b
0
;
if
(
CAHBLTlIlll
[
5
]
)
assign
CAHBLTIlI0l
=
CAHBLTlOI0l
;
else
assign
CAHBLTIlI0l
=
1
'b
0
;
if
(
CAHBLTlIlll
[
6
]
)
assign
CAHBLTlOl0l
=
CAHBLTO1I0l
;
else
assign
CAHBLTlOl0l
=
1
'b
0
;
if
(
CAHBLTlIlll
[
7
]
)
assign
CAHBLTO1l0l
=
CAHBLTIll0l
;
else
assign
CAHBLTO1l0l
=
1
'b
0
;
if
(
CAHBLTlIlll
[
8
]
)
assign
CAHBLTIl00l
=
CAHBLTlO00l
;
else
assign
CAHBLTIl00l
=
1
'b
0
;
if
(
CAHBLTlIlll
[
9
]
)
assign
CAHBLTlO10l
=
CAHBLTO100l
;
else
assign
CAHBLTlO10l
=
1
'b
0
;
if
(
CAHBLTlIlll
[
10
]
)
assign
CAHBLTO110l
=
CAHBLTIl10l
;
else
assign
CAHBLTO110l
=
1
'b
0
;
if
(
CAHBLTlIlll
[
11
]
)
assign
CAHBLTIlO1l
=
CAHBLTlOO1l
;
else
assign
CAHBLTIlO1l
=
1
'b
0
;
if
(
CAHBLTlIlll
[
12
]
)
assign
CAHBLTlOI1l
=
CAHBLTO1O1l
;
else
assign
CAHBLTlOI1l
=
1
'b
0
;
if
(
CAHBLTlIlll
[
13
]
)
assign
CAHBLTO1I1l
=
CAHBLTIlI1l
;
else
assign
CAHBLTO1I1l
=
1
'b
0
;
if
(
CAHBLTlIlll
[
14
]
)
assign
CAHBLTIll1l
=
CAHBLTlOl1l
;
else
assign
CAHBLTIll1l
=
1
'b
0
;
if
(
CAHBLTlIlll
[
15
]
)
assign
CAHBLTlO01l
=
CAHBLTO1l1l
;
else
assign
CAHBLTlO01l
=
1
'b
0
;
if
(
CAHBLTlIlll
[
16
]
)
assign
CAHBLTO101l
=
CAHBLTIl01l
;
else
assign
CAHBLTO101l
=
1
'b
0
;
if
(
CAHBLTOllll
[
0
]
)
assign
CAHBLTll11l
=
CAHBLTOI11l
;
else
assign
CAHBLTll11l
=
1
'b
0
;
if
(
CAHBLTOllll
[
1
]
)
assign
CAHBLTOIOO0
=
CAHBLTI111l
;
else
assign
CAHBLTOIOO0
=
1
'b
0
;
if
(
CAHBLTOllll
[
2
]
)
assign
CAHBLTI1OO0
=
CAHBLTllOO0
;
else
assign
CAHBLTI1OO0
=
1
'b
0
;
if
(
CAHBLTOllll
[
3
]
)
assign
CAHBLTllIO0
=
CAHBLTOIIO0
;
else
assign
CAHBLTllIO0
=
1
'b
0
;
if
(
CAHBLTOllll
[
4
]
)
assign
CAHBLTOIlO0
=
CAHBLTI1IO0
;
else
assign
CAHBLTOIlO0
=
1
'b
0
;
if
(
CAHBLTOllll
[
5
]
)
assign
CAHBLTI1lO0
=
CAHBLTlllO0
;
else
assign
CAHBLTI1lO0
=
1
'b
0
;
if
(
CAHBLTOllll
[
6
]
)
assign
CAHBLTll0O0
=
CAHBLTOI0O0
;
else
assign
CAHBLTll0O0
=
1
'b
0
;
if
(
CAHBLTOllll
[
7
]
)
assign
CAHBLTOI1O0
=
CAHBLTI10O0
;
else
assign
CAHBLTOI1O0
=
1
'b
0
;
if
(
CAHBLTOllll
[
8
]
)
assign
CAHBLTI11O0
=
CAHBLTll1O0
;
else
assign
CAHBLTI11O0
=
1
'b
0
;
if
(
CAHBLTOllll
[
9
]
)
assign
CAHBLTllOI0
=
CAHBLTOIOI0
;
else
assign
CAHBLTllOI0
=
1
'b
0
;
if
(
CAHBLTOllll
[
10
]
)
assign
CAHBLTOIII0
=
CAHBLTI1OI0
;
else
assign
CAHBLTOIII0
=
1
'b
0
;
if
(
CAHBLTOllll
[
11
]
)
assign
CAHBLTI1II0
=
CAHBLTllII0
;
else
assign
CAHBLTI1II0
=
1
'b
0
;
if
(
CAHBLTOllll
[
12
]
)
assign
CAHBLTlllI0
=
CAHBLTOIlI0
;
else
assign
CAHBLTlllI0
=
1
'b
0
;
if
(
CAHBLTOllll
[
13
]
)
assign
CAHBLTOI0I0
=
CAHBLTI1lI0
;
else
assign
CAHBLTOI0I0
=
1
'b
0
;
if
(
CAHBLTOllll
[
14
]
)
assign
CAHBLTI10I0
=
CAHBLTll0I0
;
else
assign
CAHBLTI10I0
=
1
'b
0
;
if
(
CAHBLTOllll
[
15
]
)
assign
CAHBLTll1I0
=
CAHBLTOI1I0
;
else
assign
CAHBLTll1I0
=
1
'b
0
;
if
(
CAHBLTOllll
[
16
]
)
assign
CAHBLTOIOl0
=
CAHBLTI11I0
;
else
assign
CAHBLTOIOl0
=
1
'b
0
;
endgenerate
generate
if
(
CAHBLTIIO0
[
0
]
)
assign
CAHBLTO1O0
=
CAHBLTIlO0
;
else
assign
CAHBLTO1O0
=
1
'b
0
;
if
(
CAHBLTIIO0
[
1
]
)
assign
CAHBLTIlI0
=
CAHBLTlOI0
;
else
assign
CAHBLTIlI0
=
1
'b
0
;
if
(
CAHBLTIIO0
[
2
]
)
assign
CAHBLTlOl0
=
CAHBLTO1I0
;
else
assign
CAHBLTlOl0
=
1
'b
0
;
if
(
CAHBLTIIO0
[
3
]
)
assign
CAHBLTO1l0
=
CAHBLTIll0
;
else
assign
CAHBLTO1l0
=
1
'b
0
;
if
(
CAHBLTIIO0
[
4
]
)
assign
CAHBLTIl00
=
CAHBLTlO00
;
else
assign
CAHBLTIl00
=
1
'b
0
;
if
(
CAHBLTIIO0
[
5
]
)
assign
CAHBLTlO10
=
CAHBLTO100
;
else
assign
CAHBLTlO10
=
1
'b
0
;
if
(
CAHBLTIIO0
[
6
]
)
assign
CAHBLTO110
=
CAHBLTIl10
;
else
assign
CAHBLTO110
=
1
'b
0
;
if
(
CAHBLTIIO0
[
7
]
)
assign
CAHBLTIlO1
=
CAHBLTlOO1
;
else
assign
CAHBLTIlO1
=
1
'b
0
;
if
(
CAHBLTIIO0
[
8
]
)
assign
CAHBLTlOI1
=
CAHBLTO1O1
;
else
assign
CAHBLTlOI1
=
1
'b
0
;
if
(
CAHBLTIIO0
[
9
]
)
assign
CAHBLTO1I1
=
CAHBLTIlI1
;
else
assign
CAHBLTO1I1
=
1
'b
0
;
if
(
CAHBLTIIO0
[
10
]
)
assign
CAHBLTIll1
=
CAHBLTlOl1
;
else
assign
CAHBLTIll1
=
1
'b
0
;
if
(
CAHBLTIIO0
[
11
]
)
assign
CAHBLTlO01
=
CAHBLTO1l1
;
else
assign
CAHBLTlO01
=
1
'b
0
;
if
(
CAHBLTIIO0
[
12
]
)
assign
CAHBLTO101
=
CAHBLTIl01
;
else
assign
CAHBLTO101
=
1
'b
0
;
if
(
CAHBLTIIO0
[
13
]
)
assign
CAHBLTIl11
=
CAHBLTlO11
;
else
assign
CAHBLTIl11
=
1
'b
0
;
if
(
CAHBLTIIO0
[
14
]
)
assign
CAHBLTlOOOI
=
CAHBLTO111
;
else
assign
CAHBLTlOOOI
=
1
'b
0
;
if
(
CAHBLTIIO0
[
15
]
)
assign
CAHBLTO1OOI
=
CAHBLTIlOOI
;
else
assign
CAHBLTO1OOI
=
1
'b
0
;
if
(
CAHBLTIIO0
[
16
]
)
assign
CAHBLTIlIOI
=
CAHBLTlOIOI
;
else
assign
CAHBLTIlIOI
=
1
'b
0
;
if
(
CAHBLTlIO0
[
0
]
)
assign
CAHBLTOIlOI
=
CAHBLTI1IOI
;
else
assign
CAHBLTOIlOI
=
1
'b
0
;
if
(
CAHBLTlIO0
[
1
]
)
assign
CAHBLTI1lOI
=
CAHBLTlllOI
;
else
assign
CAHBLTI1lOI
=
1
'b
0
;
if
(
CAHBLTlIO0
[
2
]
)
assign
CAHBLTll0OI
=
CAHBLTOI0OI
;
else
assign
CAHBLTll0OI
=
1
'b
0
;
if
(
CAHBLTlIO0
[
3
]
)
assign
CAHBLTOI1OI
=
CAHBLTI10OI
;
else
assign
CAHBLTOI1OI
=
1
'b
0
;
if
(
CAHBLTlIO0
[
4
]
)
assign
CAHBLTI11OI
=
CAHBLTll1OI
;
else
assign
CAHBLTI11OI
=
1
'b
0
;
if
(
CAHBLTlIO0
[
5
]
)
assign
CAHBLTllOII
=
CAHBLTOIOII
;
else
assign
CAHBLTllOII
=
1
'b
0
;
if
(
CAHBLTlIO0
[
6
]
)
assign
CAHBLTOIIII
=
CAHBLTI1OII
;
else
assign
CAHBLTOIIII
=
1
'b
0
;
if
(
CAHBLTlIO0
[
7
]
)
assign
CAHBLTI1III
=
CAHBLTllIII
;
else
assign
CAHBLTI1III
=
1
'b
0
;
if
(
CAHBLTlIO0
[
8
]
)
assign
CAHBLTlllII
=
CAHBLTOIlII
;
else
assign
CAHBLTlllII
=
1
'b
0
;
if
(
CAHBLTlIO0
[
9
]
)
assign
CAHBLTOI0II
=
CAHBLTI1lII
;
else
assign
CAHBLTOI0II
=
1
'b
0
;
if
(
CAHBLTlIO0
[
10
]
)
assign
CAHBLTI10II
=
CAHBLTll0II
;
else
assign
CAHBLTI10II
=
1
'b
0
;
if
(
CAHBLTlIO0
[
11
]
)
assign
CAHBLTll1II
=
CAHBLTOI1II
;
else
assign
CAHBLTll1II
=
1
'b
0
;
if
(
CAHBLTlIO0
[
12
]
)
assign
CAHBLTOIOlI
=
CAHBLTI11II
;
else
assign
CAHBLTOIOlI
=
1
'b
0
;
if
(
CAHBLTlIO0
[
13
]
)
assign
CAHBLTI1OlI
=
CAHBLTllOlI
;
else
assign
CAHBLTI1OlI
=
1
'b
0
;
if
(
CAHBLTlIO0
[
14
]
)
assign
CAHBLTllIlI
=
CAHBLTOIIlI
;
else
assign
CAHBLTllIlI
=
1
'b
0
;
if
(
CAHBLTlIO0
[
15
]
)
assign
CAHBLTOIllI
=
CAHBLTI1IlI
;
else
assign
CAHBLTOIllI
=
1
'b
0
;
if
(
CAHBLTlIO0
[
16
]
)
assign
CAHBLTI1llI
=
CAHBLTllllI
;
else
assign
CAHBLTI1llI
=
1
'b
0
;
if
(
CAHBLTlIlll
[
0
]
)
assign
CAHBLTI1lll
=
CAHBLTlllll
;
else
assign
CAHBLTI1lll
=
1
'b
0
;
if
(
CAHBLTlIlll
[
1
]
)
assign
CAHBLTll0ll
=
CAHBLTOI0ll
;
else
assign
CAHBLTll0ll
=
1
'b
0
;
if
(
CAHBLTlIlll
[
2
]
)
assign
CAHBLTOI1ll
=
CAHBLTI10ll
;
else
assign
CAHBLTOI1ll
=
1
'b
0
;
if
(
CAHBLTlIlll
[
3
]
)
assign
CAHBLTI11ll
=
CAHBLTll1ll
;
else
assign
CAHBLTI11ll
=
1
'b
0
;
if
(
CAHBLTlIlll
[
4
]
)
assign
CAHBLTllO0l
=
CAHBLTOIO0l
;
else
assign
CAHBLTllO0l
=
1
'b
0
;
if
(
CAHBLTlIlll
[
5
]
)
assign
CAHBLTOII0l
=
CAHBLTI1O0l
;
else
assign
CAHBLTOII0l
=
1
'b
0
;
if
(
CAHBLTlIlll
[
6
]
)
assign
CAHBLTI1I0l
=
CAHBLTllI0l
;
else
assign
CAHBLTI1I0l
=
1
'b
0
;
if
(
CAHBLTlIlll
[
7
]
)
assign
CAHBLTlll0l
=
CAHBLTOIl0l
;
else
assign
CAHBLTlll0l
=
1
'b
0
;
if
(
CAHBLTlIlll
[
8
]
)
assign
CAHBLTOI00l
=
CAHBLTI1l0l
;
else
assign
CAHBLTOI00l
=
1
'b
0
;
if
(
CAHBLTlIlll
[
9
]
)
assign
CAHBLTI100l
=
CAHBLTll00l
;
else
assign
CAHBLTI100l
=
1
'b
0
;
if
(
CAHBLTlIlll
[
10
]
)
assign
CAHBLTll10l
=
CAHBLTOI10l
;
else
assign
CAHBLTll10l
=
1
'b
0
;
if
(
CAHBLTlIlll
[
11
]
)
assign
CAHBLTOIO1l
=
CAHBLTI110l
;
else
assign
CAHBLTOIO1l
=
1
'b
0
;
if
(
CAHBLTlIlll
[
12
]
)
assign
CAHBLTI1O1l
=
CAHBLTllO1l
;
else
assign
CAHBLTI1O1l
=
1
'b
0
;
if
(
CAHBLTlIlll
[
13
]
)
assign
CAHBLTllI1l
=
CAHBLTOII1l
;
else
assign
CAHBLTllI1l
=
1
'b
0
;
if
(
CAHBLTlIlll
[
14
]
)
assign
CAHBLTOIl1l
=
CAHBLTI1I1l
;
else
assign
CAHBLTOIl1l
=
1
'b
0
;
if
(
CAHBLTlIlll
[
15
]
)
assign
CAHBLTI1l1l
=
CAHBLTlll1l
;
else
assign
CAHBLTI1l1l
=
1
'b
0
;
if
(
CAHBLTlIlll
[
16
]
)
assign
CAHBLTll01l
=
CAHBLTOI01l
;
else
assign
CAHBLTll01l
=
1
'b
0
;
if
(
CAHBLTOllll
[
0
]
)
assign
CAHBLTII11l
=
CAHBLTl101l
;
else
assign
CAHBLTII11l
=
1
'b
0
;
if
(
CAHBLTOllll
[
1
]
)
assign
CAHBLTl111l
=
CAHBLTO011l
;
else
assign
CAHBLTl111l
=
1
'b
0
;
if
(
CAHBLTOllll
[
2
]
)
assign
CAHBLTO0OO0
=
CAHBLTIIOO0
;
else
assign
CAHBLTO0OO0
=
1
'b
0
;
if
(
CAHBLTOllll
[
3
]
)
assign
CAHBLTIIIO0
=
CAHBLTl1OO0
;
else
assign
CAHBLTIIIO0
=
1
'b
0
;
if
(
CAHBLTOllll
[
4
]
)
assign
CAHBLTl1IO0
=
CAHBLTO0IO0
;
else
assign
CAHBLTl1IO0
=
1
'b
0
;
if
(
CAHBLTOllll
[
5
]
)
assign
CAHBLTO0lO0
=
CAHBLTIIlO0
;
else
assign
CAHBLTO0lO0
=
1
'b
0
;
if
(
CAHBLTOllll
[
6
]
)
assign
CAHBLTII0O0
=
CAHBLTl1lO0
;
else
assign
CAHBLTII0O0
=
1
'b
0
;
if
(
CAHBLTOllll
[
7
]
)
assign
CAHBLTl10O0
=
CAHBLTO00O0
;
else
assign
CAHBLTl10O0
=
1
'b
0
;
if
(
CAHBLTOllll
[
8
]
)
assign
CAHBLTO01O0
=
CAHBLTII1O0
;
else
assign
CAHBLTO01O0
=
1
'b
0
;
if
(
CAHBLTOllll
[
9
]
)
assign
CAHBLTIIOI0
=
CAHBLTl11O0
;
else
assign
CAHBLTIIOI0
=
1
'b
0
;
if
(
CAHBLTOllll
[
10
]
)
assign
CAHBLTl1OI0
=
CAHBLTO0OI0
;
else
assign
CAHBLTl1OI0
=
1
'b
0
;
if
(
CAHBLTOllll
[
11
]
)
assign
CAHBLTO0II0
=
CAHBLTIIII0
;
else
assign
CAHBLTO0II0
=
1
'b
0
;
if
(
CAHBLTOllll
[
12
]
)
assign
CAHBLTIIlI0
=
CAHBLTl1II0
;
else
assign
CAHBLTIIlI0
=
1
'b
0
;
if
(
CAHBLTOllll
[
13
]
)
assign
CAHBLTl1lI0
=
CAHBLTO0lI0
;
else
assign
CAHBLTl1lI0
=
1
'b
0
;
if
(
CAHBLTOllll
[
14
]
)
assign
CAHBLTO00I0
=
CAHBLTII0I0
;
else
assign
CAHBLTO00I0
=
1
'b
0
;
if
(
CAHBLTOllll
[
15
]
)
assign
CAHBLTII1I0
=
CAHBLTl10I0
;
else
assign
CAHBLTII1I0
=
1
'b
0
;
if
(
CAHBLTOllll
[
16
]
)
assign
CAHBLTl11I0
=
CAHBLTO01I0
;
else
assign
CAHBLTl11I0
=
1
'b
0
;
endgenerate
generate
if
(
CAHBLTIIO0
[
0
]
)
assign
CAHBLTI1O0
=
CAHBLTllO0
;
else
assign
CAHBLTI1O0
=
1
'b
0
;
if
(
CAHBLTIIO0
[
1
]
)
assign
CAHBLTllI0
=
CAHBLTOII0
;
else
assign
CAHBLTllI0
=
1
'b
0
;
if
(
CAHBLTIIO0
[
2
]
)
assign
CAHBLTOIl0
=
CAHBLTI1I0
;
else
assign
CAHBLTOIl0
=
1
'b
0
;
if
(
CAHBLTIIO0
[
3
]
)
assign
CAHBLTI1l0
=
CAHBLTlll0
;
else
assign
CAHBLTI1l0
=
1
'b
0
;
if
(
CAHBLTIIO0
[
4
]
)
assign
CAHBLTll00
=
CAHBLTOI00
;
else
assign
CAHBLTll00
=
1
'b
0
;
if
(
CAHBLTIIO0
[
5
]
)
assign
CAHBLTOI10
=
CAHBLTI100
;
else
assign
CAHBLTOI10
=
1
'b
0
;
if
(
CAHBLTIIO0
[
6
]
)
assign
CAHBLTI110
=
CAHBLTll10
;
else
assign
CAHBLTI110
=
1
'b
0
;
if
(
CAHBLTIIO0
[
7
]
)
assign
CAHBLTllO1
=
CAHBLTOIO1
;
else
assign
CAHBLTllO1
=
1
'b
0
;
if
(
CAHBLTIIO0
[
8
]
)
assign
CAHBLTOII1
=
CAHBLTI1O1
;
else
assign
CAHBLTOII1
=
1
'b
0
;
if
(
CAHBLTIIO0
[
9
]
)
assign
CAHBLTI1I1
=
CAHBLTllI1
;
else
assign
CAHBLTI1I1
=
1
'b
0
;
if
(
CAHBLTIIO0
[
10
]
)
assign
CAHBLTlll1
=
CAHBLTOIl1
;
else
assign
CAHBLTlll1
=
1
'b
0
;
if
(
CAHBLTIIO0
[
11
]
)
assign
CAHBLTOI01
=
CAHBLTI1l1
;
else
assign
CAHBLTOI01
=
1
'b
0
;
if
(
CAHBLTIIO0
[
12
]
)
assign
CAHBLTI101
=
CAHBLTll01
;
else
assign
CAHBLTI101
=
1
'b
0
;
if
(
CAHBLTIIO0
[
13
]
)
assign
CAHBLTll11
=
CAHBLTOI11
;
else
assign
CAHBLTll11
=
1
'b
0
;
if
(
CAHBLTIIO0
[
14
]
)
assign
CAHBLTOIOOI
=
CAHBLTI111
;
else
assign
CAHBLTOIOOI
=
1
'b
0
;
if
(
CAHBLTIIO0
[
15
]
)
assign
CAHBLTI1OOI
=
CAHBLTllOOI
;
else
assign
CAHBLTI1OOI
=
1
'b
0
;
if
(
CAHBLTIIO0
[
16
]
)
assign
CAHBLTllIOI
=
CAHBLTOIIOI
;
else
assign
CAHBLTllIOI
=
1
'b
0
;
if
(
CAHBLTlIO0
[
0
]
)
assign
CAHBLTIIlOI
=
CAHBLTl1IOI
;
else
assign
CAHBLTIIlOI
=
1
'b
0
;
if
(
CAHBLTlIO0
[
1
]
)
assign
CAHBLTl1lOI
=
CAHBLTO0lOI
;
else
assign
CAHBLTl1lOI
=
1
'b
0
;
if
(
CAHBLTlIO0
[
2
]
)
assign
CAHBLTO00OI
=
CAHBLTII0OI
;
else
assign
CAHBLTO00OI
=
1
'b
0
;
if
(
CAHBLTlIO0
[
3
]
)
assign
CAHBLTII1OI
=
CAHBLTl10OI
;
else
assign
CAHBLTII1OI
=
1
'b
0
;
if
(
CAHBLTlIO0
[
4
]
)
assign
CAHBLTl11OI
=
CAHBLTO01OI
;
else
assign
CAHBLTl11OI
=
1
'b
0
;
if
(
CAHBLTlIO0
[
5
]
)
assign
CAHBLTO0OII
=
CAHBLTIIOII
;
else
assign
CAHBLTO0OII
=
1
'b
0
;
if
(
CAHBLTlIO0
[
6
]
)
assign
CAHBLTIIIII
=
CAHBLTl1OII
;
else
assign
CAHBLTIIIII
=
1
'b
0
;
if
(
CAHBLTlIO0
[
7
]
)
assign
CAHBLTl1III
=
CAHBLTO0III
;
else
assign
CAHBLTl1III
=
1
'b
0
;
if
(
CAHBLTlIO0
[
8
]
)
assign
CAHBLTO0lII
=
CAHBLTIIlII
;
else
assign
CAHBLTO0lII
=
1
'b
0
;
if
(
CAHBLTlIO0
[
9
]
)
assign
CAHBLTII0II
=
CAHBLTl1lII
;
else
assign
CAHBLTII0II
=
1
'b
0
;
if
(
CAHBLTlIO0
[
10
]
)
assign
CAHBLTl10II
=
CAHBLTO00II
;
else
assign
CAHBLTl10II
=
1
'b
0
;
if
(
CAHBLTlIO0
[
11
]
)
assign
CAHBLTO01II
=
CAHBLTII1II
;
else
assign
CAHBLTO01II
=
1
'b
0
;
if
(
CAHBLTlIO0
[
12
]
)
assign
CAHBLTIIOlI
=
CAHBLTl11II
;
else
assign
CAHBLTIIOlI
=
1
'b
0
;
if
(
CAHBLTlIO0
[
13
]
)
assign
CAHBLTl1OlI
=
CAHBLTO0OlI
;
else
assign
CAHBLTl1OlI
=
1
'b
0
;
if
(
CAHBLTlIO0
[
14
]
)
assign
CAHBLTO0IlI
=
CAHBLTIIIlI
;
else
assign
CAHBLTO0IlI
=
1
'b
0
;
if
(
CAHBLTlIO0
[
15
]
)
assign
CAHBLTIIllI
=
CAHBLTl1IlI
;
else
assign
CAHBLTIIllI
=
1
'b
0
;
if
(
CAHBLTlIO0
[
16
]
)
assign
CAHBLTl1llI
=
CAHBLTO0llI
;
else
assign
CAHBLTl1llI
=
1
'b
0
;
if
(
CAHBLTlIlll
[
0
]
)
assign
CAHBLTl1lll
=
CAHBLTO0lll
;
else
assign
CAHBLTl1lll
=
1
'b
0
;
if
(
CAHBLTlIlll
[
1
]
)
assign
CAHBLTO00ll
=
CAHBLTII0ll
;
else
assign
CAHBLTO00ll
=
1
'b
0
;
if
(
CAHBLTlIlll
[
2
]
)
assign
CAHBLTII1ll
=
CAHBLTl10ll
;
else
assign
CAHBLTII1ll
=
1
'b
0
;
if
(
CAHBLTlIlll
[
3
]
)
assign
CAHBLTl11ll
=
CAHBLTO01ll
;
else
assign
CAHBLTl11ll
=
1
'b
0
;
if
(
CAHBLTlIlll
[
4
]
)
assign
CAHBLTO0O0l
=
CAHBLTIIO0l
;
else
assign
CAHBLTO0O0l
=
1
'b
0
;
if
(
CAHBLTlIlll
[
5
]
)
assign
CAHBLTIII0l
=
CAHBLTl1O0l
;
else
assign
CAHBLTIII0l
=
1
'b
0
;
if
(
CAHBLTlIlll
[
6
]
)
assign
CAHBLTl1I0l
=
CAHBLTO0I0l
;
else
assign
CAHBLTl1I0l
=
1
'b
0
;
if
(
CAHBLTlIlll
[
7
]
)
assign
CAHBLTO0l0l
=
CAHBLTIIl0l
;
else
assign
CAHBLTO0l0l
=
1
'b
0
;
if
(
CAHBLTlIlll
[
8
]
)
assign
CAHBLTII00l
=
CAHBLTl1l0l
;
else
assign
CAHBLTII00l
=
1
'b
0
;
if
(
CAHBLTlIlll
[
9
]
)
assign
CAHBLTl100l
=
CAHBLTO000l
;
else
assign
CAHBLTl100l
=
1
'b
0
;
if
(
CAHBLTlIlll
[
10
]
)
assign
CAHBLTO010l
=
CAHBLTII10l
;
else
assign
CAHBLTO010l
=
1
'b
0
;
if
(
CAHBLTlIlll
[
11
]
)
assign
CAHBLTIIO1l
=
CAHBLTl110l
;
else
assign
CAHBLTIIO1l
=
1
'b
0
;
if
(
CAHBLTlIlll
[
12
]
)
assign
CAHBLTl1O1l
=
CAHBLTO0O1l
;
else
assign
CAHBLTl1O1l
=
1
'b
0
;
if
(
CAHBLTlIlll
[
13
]
)
assign
CAHBLTO0I1l
=
CAHBLTIII1l
;
else
assign
CAHBLTO0I1l
=
1
'b
0
;
if
(
CAHBLTlIlll
[
14
]
)
assign
CAHBLTIIl1l
=
CAHBLTl1I1l
;
else
assign
CAHBLTIIl1l
=
1
'b
0
;
if
(
CAHBLTlIlll
[
15
]
)
assign
CAHBLTl1l1l
=
CAHBLTO0l1l
;
else
assign
CAHBLTl1l1l
=
1
'b
0
;
if
(
CAHBLTlIlll
[
16
]
)
assign
CAHBLTO001l
=
CAHBLTII01l
;
else
assign
CAHBLTO001l
=
1
'b
0
;
if
(
CAHBLTOllll
[
0
]
)
assign
CAHBLTlI11l
=
CAHBLTOO11l
;
else
assign
CAHBLTlI11l
=
1
'b
0
;
if
(
CAHBLTOllll
[
1
]
)
assign
CAHBLTOOOO0
=
CAHBLTI011l
;
else
assign
CAHBLTOOOO0
=
1
'b
0
;
if
(
CAHBLTOllll
[
2
]
)
assign
CAHBLTI0OO0
=
CAHBLTlIOO0
;
else
assign
CAHBLTI0OO0
=
1
'b
0
;
if
(
CAHBLTOllll
[
3
]
)
assign
CAHBLTlIIO0
=
CAHBLTOOIO0
;
else
assign
CAHBLTlIIO0
=
1
'b
0
;
if
(
CAHBLTOllll
[
4
]
)
assign
CAHBLTOOlO0
=
CAHBLTI0IO0
;
else
assign
CAHBLTOOlO0
=
1
'b
0
;
if
(
CAHBLTOllll
[
5
]
)
assign
CAHBLTI0lO0
=
CAHBLTlIlO0
;
else
assign
CAHBLTI0lO0
=
1
'b
0
;
if
(
CAHBLTOllll
[
6
]
)
assign
CAHBLTlI0O0
=
CAHBLTOO0O0
;
else
assign
CAHBLTlI0O0
=
1
'b
0
;
if
(
CAHBLTOllll
[
7
]
)
assign
CAHBLTOO1O0
=
CAHBLTI00O0
;
else
assign
CAHBLTOO1O0
=
1
'b
0
;
if
(
CAHBLTOllll
[
8
]
)
assign
CAHBLTI01O0
=
CAHBLTlI1O0
;
else
assign
CAHBLTI01O0
=
1
'b
0
;
if
(
CAHBLTOllll
[
9
]
)
assign
CAHBLTlIOI0
=
CAHBLTOOOI0
;
else
assign
CAHBLTlIOI0
=
1
'b
0
;
if
(
CAHBLTOllll
[
10
]
)
assign
CAHBLTOOII0
=
CAHBLTI0OI0
;
else
assign
CAHBLTOOII0
=
1
'b
0
;
if
(
CAHBLTOllll
[
11
]
)
assign
CAHBLTI0II0
=
CAHBLTlIII0
;
else
assign
CAHBLTI0II0
=
1
'b
0
;
if
(
CAHBLTOllll
[
12
]
)
assign
CAHBLTlIlI0
=
CAHBLTOOlI0
;
else
assign
CAHBLTlIlI0
=
1
'b
0
;
if
(
CAHBLTOllll
[
13
]
)
assign
CAHBLTOO0I0
=
CAHBLTI0lI0
;
else
assign
CAHBLTOO0I0
=
1
'b
0
;
if
(
CAHBLTOllll
[
14
]
)
assign
CAHBLTI00I0
=
CAHBLTlI0I0
;
else
assign
CAHBLTI00I0
=
1
'b
0
;
if
(
CAHBLTOllll
[
15
]
)
assign
CAHBLTlI1I0
=
CAHBLTOO1I0
;
else
assign
CAHBLTlI1I0
=
1
'b
0
;
if
(
CAHBLTOllll
[
16
]
)
assign
CAHBLTOOOl0
=
CAHBLTI01I0
;
else
assign
CAHBLTOOOl0
=
1
'b
0
;
endgenerate
generate
if
(
CAHBLTIIO0
[
0
]
)
assign
CAHBLTIIl1I
=
CAHBLTI11I
;
else
assign
CAHBLTIIl1I
=
32
'h
0
;
if
(
CAHBLTIIO0
[
1
]
)
assign
CAHBLTlIl1I
=
CAHBLTI11I
;
else
assign
CAHBLTlIl1I
=
32
'h
0
;
if
(
CAHBLTIIO0
[
2
]
)
assign
CAHBLTOll1I
=
CAHBLTI11I
;
else
assign
CAHBLTOll1I
=
32
'h
0
;
if
(
CAHBLTIIO0
[
3
]
)
assign
CAHBLTIll1I
=
CAHBLTI11I
;
else
assign
CAHBLTIll1I
=
32
'h
0
;
if
(
CAHBLTIIO0
[
4
]
)
assign
CAHBLTlll1I
=
CAHBLTI11I
;
else
assign
CAHBLTlll1I
=
32
'h
0
;
if
(
CAHBLTIIO0
[
5
]
)
assign
CAHBLTO0l1I
=
CAHBLTI11I
;
else
assign
CAHBLTO0l1I
=
32
'h
0
;
if
(
CAHBLTIIO0
[
6
]
)
assign
CAHBLTI0l1I
=
CAHBLTI11I
;
else
assign
CAHBLTI0l1I
=
32
'h
0
;
if
(
CAHBLTIIO0
[
7
]
)
assign
CAHBLTl0l1I
=
CAHBLTI11I
;
else
assign
CAHBLTl0l1I
=
32
'h
0
;
if
(
CAHBLTIIO0
[
8
]
)
assign
CAHBLTO1l1I
=
CAHBLTI11I
;
else
assign
CAHBLTO1l1I
=
32
'h
0
;
if
(
CAHBLTIIO0
[
9
]
)
assign
CAHBLTI1l1I
=
CAHBLTI11I
;
else
assign
CAHBLTI1l1I
=
32
'h
0
;
if
(
CAHBLTIIO0
[
10
]
)
assign
CAHBLTl1l1I
=
CAHBLTI11I
;
else
assign
CAHBLTl1l1I
=
32
'h
0
;
if
(
CAHBLTIIO0
[
11
]
)
assign
CAHBLTOO01I
=
CAHBLTI11I
;
else
assign
CAHBLTOO01I
=
32
'h
0
;
if
(
CAHBLTIIO0
[
12
]
)
assign
CAHBLTIO01I
=
CAHBLTI11I
;
else
assign
CAHBLTIO01I
=
32
'h
0
;
if
(
CAHBLTIIO0
[
13
]
)
assign
CAHBLTlO01I
=
CAHBLTI11I
;
else
assign
CAHBLTlO01I
=
32
'h
0
;
if
(
CAHBLTIIO0
[
14
]
)
assign
CAHBLTOI01I
=
CAHBLTI11I
;
else
assign
CAHBLTOI01I
=
32
'h
0
;
if
(
CAHBLTIIO0
[
15
]
)
assign
CAHBLTII01I
=
CAHBLTI11I
;
else
assign
CAHBLTII01I
=
32
'h
0
;
if
(
CAHBLTIIO0
[
16
]
)
assign
CAHBLTlI01I
=
CAHBLTI11I
;
else
assign
CAHBLTlI01I
=
32
'h
0
;
if
(
CAHBLTlIO0
[
0
]
)
assign
CAHBLTOl01I
=
CAHBLTlOOl
;
else
assign
CAHBLTOl01I
=
32
'h
0
;
if
(
CAHBLTlIO0
[
1
]
)
assign
CAHBLTIl01I
=
CAHBLTlOOl
;
else
assign
CAHBLTIl01I
=
32
'h
0
;
if
(
CAHBLTlIO0
[
2
]
)
assign
CAHBLTll01I
=
CAHBLTlOOl
;
else
assign
CAHBLTll01I
=
32
'h
0
;
if
(
CAHBLTlIO0
[
3
]
)
assign
CAHBLTO001I
=
CAHBLTlOOl
;
else
assign
CAHBLTO001I
=
32
'h
0
;
if
(
CAHBLTlIO0
[
4
]
)
assign
CAHBLTI001I
=
CAHBLTlOOl
;
else
assign
CAHBLTI001I
=
32
'h
0
;
if
(
CAHBLTlIO0
[
5
]
)
assign
CAHBLTl001I
=
CAHBLTlOOl
;
else
assign
CAHBLTl001I
=
32
'h
0
;
if
(
CAHBLTlIO0
[
6
]
)
assign
CAHBLTO101I
=
CAHBLTlOOl
;
else
assign
CAHBLTO101I
=
32
'h
0
;
if
(
CAHBLTlIO0
[
7
]
)
assign
CAHBLTI101I
=
CAHBLTlOOl
;
else
assign
CAHBLTI101I
=
32
'h
0
;
if
(
CAHBLTlIO0
[
8
]
)
assign
CAHBLTl101I
=
CAHBLTlOOl
;
else
assign
CAHBLTl101I
=
32
'h
0
;
if
(
CAHBLTlIO0
[
9
]
)
assign
CAHBLTOO11I
=
CAHBLTlOOl
;
else
assign
CAHBLTOO11I
=
32
'h
0
;
if
(
CAHBLTlIO0
[
10
]
)
assign
CAHBLTIO11I
=
CAHBLTlOOl
;
else
assign
CAHBLTIO11I
=
32
'h
0
;
if
(
CAHBLTlIO0
[
11
]
)
assign
CAHBLTlO11I
=
CAHBLTlOOl
;
else
assign
CAHBLTlO11I
=
32
'h
0
;
if
(
CAHBLTlIO0
[
12
]
)
assign
CAHBLTOI11I
=
CAHBLTlOOl
;
else
assign
CAHBLTOI11I
=
32
'h
0
;
if
(
CAHBLTlIO0
[
13
]
)
assign
CAHBLTII11I
=
CAHBLTlOOl
;
else
assign
CAHBLTII11I
=
32
'h
0
;
if
(
CAHBLTlIO0
[
14
]
)
assign
CAHBLTlI11I
=
CAHBLTlOOl
;
else
assign
CAHBLTlI11I
=
32
'h
0
;
if
(
CAHBLTlIO0
[
15
]
)
assign
CAHBLTOl11I
=
CAHBLTlOOl
;
else
assign
CAHBLTOl11I
=
32
'h
0
;
if
(
CAHBLTlIO0
[
16
]
)
assign
CAHBLTIl11I
=
CAHBLTlOOl
;
else
assign
CAHBLTIl11I
=
32
'h
0
;
if
(
CAHBLTlIlll
[
0
]
)
assign
CAHBLTIOl00
=
CAHBLTOlOl
;
else
assign
CAHBLTIOl00
=
32
'h
0
;
if
(
CAHBLTlIlll
[
1
]
)
assign
CAHBLTlOl00
=
CAHBLTOlOl
;
else
assign
CAHBLTlOl00
=
32
'h
0
;
if
(
CAHBLTlIlll
[
2
]
)
assign
CAHBLTOIl00
=
CAHBLTOlOl
;
else
assign
CAHBLTOIl00
=
32
'h
0
;
if
(
CAHBLTlIlll
[
3
]
)
assign
CAHBLTIIl00
=
CAHBLTOlOl
;
else
assign
CAHBLTIIl00
=
32
'h
0
;
if
(
CAHBLTlIlll
[
4
]
)
assign
CAHBLTlIl00
=
CAHBLTOlOl
;
else
assign
CAHBLTlIl00
=
32
'h
0
;
if
(
CAHBLTlIlll
[
5
]
)
assign
CAHBLTOll00
=
CAHBLTOlOl
;
else
assign
CAHBLTOll00
=
32
'h
0
;
if
(
CAHBLTlIlll
[
6
]
)
assign
CAHBLTIll00
=
CAHBLTOlOl
;
else
assign
CAHBLTIll00
=
32
'h
0
;
if
(
CAHBLTlIlll
[
7
]
)
assign
CAHBLTlll00
=
CAHBLTOlOl
;
else
assign
CAHBLTlll00
=
32
'h
0
;
if
(
CAHBLTlIlll
[
8
]
)
assign
CAHBLTO0l00
=
CAHBLTOlOl
;
else
assign
CAHBLTO0l00
=
32
'h
0
;
if
(
CAHBLTlIlll
[
9
]
)
assign
CAHBLTI0l00
=
CAHBLTOlOl
;
else
assign
CAHBLTI0l00
=
32
'h
0
;
if
(
CAHBLTlIlll
[
10
]
)
assign
CAHBLTl0l00
=
CAHBLTOlOl
;
else
assign
CAHBLTl0l00
=
32
'h
0
;
if
(
CAHBLTlIlll
[
11
]
)
assign
CAHBLTO1l00
=
CAHBLTOlOl
;
else
assign
CAHBLTO1l00
=
32
'h
0
;
if
(
CAHBLTlIlll
[
12
]
)
assign
CAHBLTI1l00
=
CAHBLTOlOl
;
else
assign
CAHBLTI1l00
=
32
'h
0
;
if
(
CAHBLTlIlll
[
13
]
)
assign
CAHBLTl1l00
=
CAHBLTOlOl
;
else
assign
CAHBLTl1l00
=
32
'h
0
;
if
(
CAHBLTlIlll
[
14
]
)
assign
CAHBLTOO000
=
CAHBLTOlOl
;
else
assign
CAHBLTOO000
=
32
'h
0
;
if
(
CAHBLTlIlll
[
15
]
)
assign
CAHBLTIO000
=
CAHBLTOlOl
;
else
assign
CAHBLTIO000
=
32
'h
0
;
if
(
CAHBLTlIlll
[
16
]
)
assign
CAHBLTlO000
=
CAHBLTOlOl
;
else
assign
CAHBLTlO000
=
32
'h
0
;
if
(
CAHBLTOllll
[
0
]
)
assign
CAHBLTOI000
=
CAHBLTI0Ol
;
else
assign
CAHBLTOI000
=
32
'h
0
;
if
(
CAHBLTOllll
[
1
]
)
assign
CAHBLTII000
=
CAHBLTI0Ol
;
else
assign
CAHBLTII000
=
32
'h
0
;
if
(
CAHBLTOllll
[
2
]
)
assign
CAHBLTlI000
=
CAHBLTI0Ol
;
else
assign
CAHBLTlI000
=
32
'h
0
;
if
(
CAHBLTOllll
[
3
]
)
assign
CAHBLTOl000
=
CAHBLTI0Ol
;
else
assign
CAHBLTOl000
=
32
'h
0
;
if
(
CAHBLTOllll
[
4
]
)
assign
CAHBLTIl000
=
CAHBLTI0Ol
;
else
assign
CAHBLTIl000
=
32
'h
0
;
if
(
CAHBLTOllll
[
5
]
)
assign
CAHBLTll000
=
CAHBLTI0Ol
;
else
assign
CAHBLTll000
=
32
'h
0
;
if
(
CAHBLTOllll
[
6
]
)
assign
CAHBLTO0000
=
CAHBLTI0Ol
;
else
assign
CAHBLTO0000
=
32
'h
0
;
if
(
CAHBLTOllll
[
7
]
)
assign
CAHBLTI0000
=
CAHBLTI0Ol
;
else
assign
CAHBLTI0000
=
32
'h
0
;
if
(
CAHBLTOllll
[
8
]
)
assign
CAHBLTl0000
=
CAHBLTI0Ol
;
else
assign
CAHBLTl0000
=
32
'h
0
;
if
(
CAHBLTOllll
[
9
]
)
assign
CAHBLTO1000
=
CAHBLTI0Ol
;
else
assign
CAHBLTO1000
=
32
'h
0
;
if
(
CAHBLTOllll
[
10
]
)
assign
CAHBLTI1000
=
CAHBLTI0Ol
;
else
assign
CAHBLTI1000
=
32
'h
0
;
if
(
CAHBLTOllll
[
11
]
)
assign
CAHBLTl1000
=
CAHBLTI0Ol
;
else
assign
CAHBLTl1000
=
32
'h
0
;
if
(
CAHBLTOllll
[
12
]
)
assign
CAHBLTOO100
=
CAHBLTI0Ol
;
else
assign
CAHBLTOO100
=
32
'h
0
;
if
(
CAHBLTOllll
[
13
]
)
assign
CAHBLTIO100
=
CAHBLTI0Ol
;
else
assign
CAHBLTIO100
=
32
'h
0
;
if
(
CAHBLTOllll
[
14
]
)
assign
CAHBLTlO100
=
CAHBLTI0Ol
;
else
assign
CAHBLTlO100
=
32
'h
0
;
if
(
CAHBLTOllll
[
15
]
)
assign
CAHBLTOI100
=
CAHBLTI0Ol
;
else
assign
CAHBLTOI100
=
32
'h
0
;
if
(
CAHBLTOllll
[
16
]
)
assign
CAHBLTII100
=
CAHBLTI0Ol
;
else
assign
CAHBLTII100
=
32
'h
0
;
endgenerate
generate
if
(
CAHBLTIIO0
[
0
]
)
assign
CAHBLTO1IOl
=
CAHBLTlI0
;
else
assign
CAHBLTO1IOl
=
1
'b
0
;
if
(
CAHBLTIIO0
[
1
]
)
assign
CAHBLTI1IOl
=
CAHBLTlI0
;
else
assign
CAHBLTI1IOl
=
1
'b
0
;
if
(
CAHBLTIIO0
[
2
]
)
assign
CAHBLTl1IOl
=
CAHBLTlI0
;
else
assign
CAHBLTl1IOl
=
1
'b
0
;
if
(
CAHBLTIIO0
[
3
]
)
assign
CAHBLTOOlOl
=
CAHBLTlI0
;
else
assign
CAHBLTOOlOl
=
1
'b
0
;
if
(
CAHBLTIIO0
[
4
]
)
assign
CAHBLTIOlOl
=
CAHBLTlI0
;
else
assign
CAHBLTIOlOl
=
1
'b
0
;
if
(
CAHBLTIIO0
[
5
]
)
assign
CAHBLTlOlOl
=
CAHBLTlI0
;
else
assign
CAHBLTlOlOl
=
1
'b
0
;
if
(
CAHBLTIIO0
[
6
]
)
assign
CAHBLTOIlOl
=
CAHBLTlI0
;
else
assign
CAHBLTOIlOl
=
1
'b
0
;
if
(
CAHBLTIIO0
[
7
]
)
assign
CAHBLTIIlOl
=
CAHBLTlI0
;
else
assign
CAHBLTIIlOl
=
1
'b
0
;
if
(
CAHBLTIIO0
[
8
]
)
assign
CAHBLTlIlOl
=
CAHBLTlI0
;
else
assign
CAHBLTlIlOl
=
1
'b
0
;
if
(
CAHBLTIIO0
[
9
]
)
assign
CAHBLTOllOl
=
CAHBLTlI0
;
else
assign
CAHBLTOllOl
=
1
'b
0
;
if
(
CAHBLTIIO0
[
10
]
)
assign
CAHBLTIllOl
=
CAHBLTlI0
;
else
assign
CAHBLTIllOl
=
1
'b
0
;
if
(
CAHBLTIIO0
[
11
]
)
assign
CAHBLTlllOl
=
CAHBLTlI0
;
else
assign
CAHBLTlllOl
=
1
'b
0
;
if
(
CAHBLTIIO0
[
12
]
)
assign
CAHBLTO0lOl
=
CAHBLTlI0
;
else
assign
CAHBLTO0lOl
=
1
'b
0
;
if
(
CAHBLTIIO0
[
13
]
)
assign
CAHBLTI0lOl
=
CAHBLTlI0
;
else
assign
CAHBLTI0lOl
=
1
'b
0
;
if
(
CAHBLTIIO0
[
14
]
)
assign
CAHBLTl0lOl
=
CAHBLTlI0
;
else
assign
CAHBLTl0lOl
=
1
'b
0
;
if
(
CAHBLTIIO0
[
15
]
)
assign
CAHBLTO1lOl
=
CAHBLTlI0
;
else
assign
CAHBLTO1lOl
=
1
'b
0
;
if
(
CAHBLTIIO0
[
16
]
)
assign
CAHBLTI1lOl
=
CAHBLTlI0
;
else
assign
CAHBLTI1lOl
=
1
'b
0
;
if
(
CAHBLTlIO0
[
0
]
)
assign
CAHBLTl1lOl
=
CAHBLTOl0
;
else
assign
CAHBLTl1lOl
=
1
'b
0
;
if
(
CAHBLTlIO0
[
1
]
)
assign
CAHBLTOO0Ol
=
CAHBLTOl0
;
else
assign
CAHBLTOO0Ol
=
1
'b
0
;
if
(
CAHBLTlIO0
[
2
]
)
assign
CAHBLTIO0Ol
=
CAHBLTOl0
;
else
assign
CAHBLTIO0Ol
=
1
'b
0
;
if
(
CAHBLTlIO0
[
3
]
)
assign
CAHBLTlO0Ol
=
CAHBLTOl0
;
else
assign
CAHBLTlO0Ol
=
1
'b
0
;
if
(
CAHBLTlIO0
[
4
]
)
assign
CAHBLTOI0Ol
=
CAHBLTOl0
;
else
assign
CAHBLTOI0Ol
=
1
'b
0
;
if
(
CAHBLTlIO0
[
5
]
)
assign
CAHBLTII0Ol
=
CAHBLTOl0
;
else
assign
CAHBLTII0Ol
=
1
'b
0
;
if
(
CAHBLTlIO0
[
6
]
)
assign
CAHBLTlI0Ol
=
CAHBLTOl0
;
else
assign
CAHBLTlI0Ol
=
1
'b
0
;
if
(
CAHBLTlIO0
[
7
]
)
assign
CAHBLTOl0Ol
=
CAHBLTOl0
;
else
assign
CAHBLTOl0Ol
=
1
'b
0
;
if
(
CAHBLTlIO0
[
8
]
)
assign
CAHBLTIl0Ol
=
CAHBLTOl0
;
else
assign
CAHBLTIl0Ol
=
1
'b
0
;
if
(
CAHBLTlIO0
[
9
]
)
assign
CAHBLTll0Ol
=
CAHBLTOl0
;
else
assign
CAHBLTll0Ol
=
1
'b
0
;
if
(
CAHBLTlIO0
[
10
]
)
assign
CAHBLTO00Ol
=
CAHBLTOl0
;
else
assign
CAHBLTO00Ol
=
1
'b
0
;
if
(
CAHBLTlIO0
[
11
]
)
assign
CAHBLTI00Ol
=
CAHBLTOl0
;
else
assign
CAHBLTI00Ol
=
1
'b
0
;
if
(
CAHBLTlIO0
[
12
]
)
assign
CAHBLTl00Ol
=
CAHBLTOl0
;
else
assign
CAHBLTl00Ol
=
1
'b
0
;
if
(
CAHBLTlIO0
[
13
]
)
assign
CAHBLTO10Ol
=
CAHBLTOl0
;
else
assign
CAHBLTO10Ol
=
1
'b
0
;
if
(
CAHBLTlIO0
[
14
]
)
assign
CAHBLTI10Ol
=
CAHBLTOl0
;
else
assign
CAHBLTI10Ol
=
1
'b
0
;
if
(
CAHBLTlIO0
[
15
]
)
assign
CAHBLTl10Ol
=
CAHBLTOl0
;
else
assign
CAHBLTl10Ol
=
1
'b
0
;
if
(
CAHBLTlIO0
[
16
]
)
assign
CAHBLTOO1Ol
=
CAHBLTOl0
;
else
assign
CAHBLTOO1Ol
=
1
'b
0
;
if
(
CAHBLTlIlll
[
0
]
)
assign
CAHBLTO0I10
=
CAHBLTIl0
;
else
assign
CAHBLTO0I10
=
1
'b
0
;
if
(
CAHBLTlIlll
[
1
]
)
assign
CAHBLTI0I10
=
CAHBLTIl0
;
else
assign
CAHBLTI0I10
=
1
'b
0
;
if
(
CAHBLTlIlll
[
2
]
)
assign
CAHBLTl0I10
=
CAHBLTIl0
;
else
assign
CAHBLTl0I10
=
1
'b
0
;
if
(
CAHBLTlIlll
[
3
]
)
assign
CAHBLTO1I10
=
CAHBLTIl0
;
else
assign
CAHBLTO1I10
=
1
'b
0
;
if
(
CAHBLTlIlll
[
4
]
)
assign
CAHBLTI1I10
=
CAHBLTIl0
;
else
assign
CAHBLTI1I10
=
1
'b
0
;
if
(
CAHBLTlIlll
[
5
]
)
assign
CAHBLTl1I10
=
CAHBLTIl0
;
else
assign
CAHBLTl1I10
=
1
'b
0
;
if
(
CAHBLTlIlll
[
6
]
)
assign
CAHBLTOOl10
=
CAHBLTIl0
;
else
assign
CAHBLTOOl10
=
1
'b
0
;
if
(
CAHBLTlIlll
[
7
]
)
assign
CAHBLTIOl10
=
CAHBLTIl0
;
else
assign
CAHBLTIOl10
=
1
'b
0
;
if
(
CAHBLTlIlll
[
8
]
)
assign
CAHBLTlOl10
=
CAHBLTIl0
;
else
assign
CAHBLTlOl10
=
1
'b
0
;
if
(
CAHBLTlIlll
[
9
]
)
assign
CAHBLTOIl10
=
CAHBLTIl0
;
else
assign
CAHBLTOIl10
=
1
'b
0
;
if
(
CAHBLTlIlll
[
10
]
)
assign
CAHBLTIIl10
=
CAHBLTIl0
;
else
assign
CAHBLTIIl10
=
1
'b
0
;
if
(
CAHBLTlIlll
[
11
]
)
assign
CAHBLTlIl10
=
CAHBLTIl0
;
else
assign
CAHBLTlIl10
=
1
'b
0
;
if
(
CAHBLTlIlll
[
12
]
)
assign
CAHBLTOll10
=
CAHBLTIl0
;
else
assign
CAHBLTOll10
=
1
'b
0
;
if
(
CAHBLTlIlll
[
13
]
)
assign
CAHBLTIll10
=
CAHBLTIl0
;
else
assign
CAHBLTIll10
=
1
'b
0
;
if
(
CAHBLTlIlll
[
14
]
)
assign
CAHBLTlll10
=
CAHBLTIl0
;
else
assign
CAHBLTlll10
=
1
'b
0
;
if
(
CAHBLTlIlll
[
15
]
)
assign
CAHBLTO0l10
=
CAHBLTIl0
;
else
assign
CAHBLTO0l10
=
1
'b
0
;
if
(
CAHBLTlIlll
[
16
]
)
assign
CAHBLTI0l10
=
CAHBLTIl0
;
else
assign
CAHBLTI0l10
=
1
'b
0
;
if
(
CAHBLTOllll
[
0
]
)
assign
CAHBLTl0l10
=
CAHBLTll0
;
else
assign
CAHBLTl0l10
=
1
'b
0
;
if
(
CAHBLTOllll
[
1
]
)
assign
CAHBLTO1l10
=
CAHBLTll0
;
else
assign
CAHBLTO1l10
=
1
'b
0
;
if
(
CAHBLTOllll
[
2
]
)
assign
CAHBLTI1l10
=
CAHBLTll0
;
else
assign
CAHBLTI1l10
=
1
'b
0
;
if
(
CAHBLTOllll
[
3
]
)
assign
CAHBLTl1l10
=
CAHBLTll0
;
else
assign
CAHBLTl1l10
=
1
'b
0
;
if
(
CAHBLTOllll
[
4
]
)
assign
CAHBLTOO010
=
CAHBLTll0
;
else
assign
CAHBLTOO010
=
1
'b
0
;
if
(
CAHBLTOllll
[
5
]
)
assign
CAHBLTIO010
=
CAHBLTll0
;
else
assign
CAHBLTIO010
=
1
'b
0
;
if
(
CAHBLTOllll
[
6
]
)
assign
CAHBLTlO010
=
CAHBLTll0
;
else
assign
CAHBLTlO010
=
1
'b
0
;
if
(
CAHBLTOllll
[
7
]
)
assign
CAHBLTOI010
=
CAHBLTll0
;
else
assign
CAHBLTOI010
=
1
'b
0
;
if
(
CAHBLTOllll
[
8
]
)
assign
CAHBLTII010
=
CAHBLTll0
;
else
assign
CAHBLTII010
=
1
'b
0
;
if
(
CAHBLTOllll
[
9
]
)
assign
CAHBLTlI010
=
CAHBLTll0
;
else
assign
CAHBLTlI010
=
1
'b
0
;
if
(
CAHBLTOllll
[
10
]
)
assign
CAHBLTOl010
=
CAHBLTll0
;
else
assign
CAHBLTOl010
=
1
'b
0
;
if
(
CAHBLTOllll
[
11
]
)
assign
CAHBLTIl010
=
CAHBLTll0
;
else
assign
CAHBLTIl010
=
1
'b
0
;
if
(
CAHBLTOllll
[
12
]
)
assign
CAHBLTll010
=
CAHBLTll0
;
else
assign
CAHBLTll010
=
1
'b
0
;
if
(
CAHBLTOllll
[
13
]
)
assign
CAHBLTO0010
=
CAHBLTll0
;
else
assign
CAHBLTO0010
=
1
'b
0
;
if
(
CAHBLTOllll
[
14
]
)
assign
CAHBLTI0010
=
CAHBLTll0
;
else
assign
CAHBLTI0010
=
1
'b
0
;
if
(
CAHBLTOllll
[
15
]
)
assign
CAHBLTl0010
=
CAHBLTll0
;
else
assign
CAHBLTl0010
=
1
'b
0
;
if
(
CAHBLTOllll
[
16
]
)
assign
CAHBLTO1010
=
CAHBLTll0
;
else
assign
CAHBLTO1010
=
1
'b
0
;
endgenerate
generate
if
(
CAHBLTIIO0
[
0
]
)
assign
CAHBLTll11I
=
CAHBLTl11I
;
else
assign
CAHBLTll11I
=
1
'b
0
;
if
(
CAHBLTIIO0
[
1
]
)
assign
CAHBLTO011I
=
CAHBLTl11I
;
else
assign
CAHBLTO011I
=
1
'b
0
;
if
(
CAHBLTIIO0
[
2
]
)
assign
CAHBLTI011I
=
CAHBLTl11I
;
else
assign
CAHBLTI011I
=
1
'b
0
;
if
(
CAHBLTIIO0
[
3
]
)
assign
CAHBLTl011I
=
CAHBLTl11I
;
else
assign
CAHBLTl011I
=
1
'b
0
;
if
(
CAHBLTIIO0
[
4
]
)
assign
CAHBLTO111I
=
CAHBLTl11I
;
else
assign
CAHBLTO111I
=
1
'b
0
;
if
(
CAHBLTIIO0
[
5
]
)
assign
CAHBLTI111I
=
CAHBLTl11I
;
else
assign
CAHBLTI111I
=
1
'b
0
;
if
(
CAHBLTIIO0
[
6
]
)
assign
CAHBLTl111I
=
CAHBLTl11I
;
else
assign
CAHBLTl111I
=
1
'b
0
;
if
(
CAHBLTIIO0
[
7
]
)
assign
CAHBLTOOOOl
=
CAHBLTl11I
;
else
assign
CAHBLTOOOOl
=
1
'b
0
;
if
(
CAHBLTIIO0
[
8
]
)
assign
CAHBLTIOOOl
=
CAHBLTl11I
;
else
assign
CAHBLTIOOOl
=
1
'b
0
;
if
(
CAHBLTIIO0
[
9
]
)
assign
CAHBLTlOOOl
=
CAHBLTl11I
;
else
assign
CAHBLTlOOOl
=
1
'b
0
;
if
(
CAHBLTIIO0
[
10
]
)
assign
CAHBLTOIOOl
=
CAHBLTl11I
;
else
assign
CAHBLTOIOOl
=
1
'b
0
;
if
(
CAHBLTIIO0
[
11
]
)
assign
CAHBLTIIOOl
=
CAHBLTl11I
;
else
assign
CAHBLTIIOOl
=
1
'b
0
;
if
(
CAHBLTIIO0
[
12
]
)
assign
CAHBLTlIOOl
=
CAHBLTl11I
;
else
assign
CAHBLTlIOOl
=
1
'b
0
;
if
(
CAHBLTIIO0
[
13
]
)
assign
CAHBLTOlOOl
=
CAHBLTl11I
;
else
assign
CAHBLTOlOOl
=
1
'b
0
;
if
(
CAHBLTIIO0
[
14
]
)
assign
CAHBLTIlOOl
=
CAHBLTl11I
;
else
assign
CAHBLTIlOOl
=
1
'b
0
;
if
(
CAHBLTIIO0
[
15
]
)
assign
CAHBLTllOOl
=
CAHBLTl11I
;
else
assign
CAHBLTllOOl
=
1
'b
0
;
if
(
CAHBLTIIO0
[
16
]
)
assign
CAHBLTO0OOl
=
CAHBLTl11I
;
else
assign
CAHBLTO0OOl
=
1
'b
0
;
if
(
CAHBLTlIO0
[
0
]
)
assign
CAHBLTI0OOl
=
CAHBLTOIOl
;
else
assign
CAHBLTI0OOl
=
1
'b
0
;
if
(
CAHBLTlIO0
[
1
]
)
assign
CAHBLTl0OOl
=
CAHBLTOIOl
;
else
assign
CAHBLTl0OOl
=
1
'b
0
;
if
(
CAHBLTlIO0
[
2
]
)
assign
CAHBLTO1OOl
=
CAHBLTOIOl
;
else
assign
CAHBLTO1OOl
=
1
'b
0
;
if
(
CAHBLTlIO0
[
3
]
)
assign
CAHBLTI1OOl
=
CAHBLTOIOl
;
else
assign
CAHBLTI1OOl
=
1
'b
0
;
if
(
CAHBLTlIO0
[
4
]
)
assign
CAHBLTl1OOl
=
CAHBLTOIOl
;
else
assign
CAHBLTl1OOl
=
1
'b
0
;
if
(
CAHBLTlIO0
[
5
]
)
assign
CAHBLTOOIOl
=
CAHBLTOIOl
;
else
assign
CAHBLTOOIOl
=
1
'b
0
;
if
(
CAHBLTlIO0
[
6
]
)
assign
CAHBLTIOIOl
=
CAHBLTOIOl
;
else
assign
CAHBLTIOIOl
=
1
'b
0
;
if
(
CAHBLTlIO0
[
7
]
)
assign
CAHBLTlOIOl
=
CAHBLTOIOl
;
else
assign
CAHBLTlOIOl
=
1
'b
0
;
if
(
CAHBLTlIO0
[
8
]
)
assign
CAHBLTOIIOl
=
CAHBLTOIOl
;
else
assign
CAHBLTOIIOl
=
1
'b
0
;
if
(
CAHBLTlIO0
[
9
]
)
assign
CAHBLTIIIOl
=
CAHBLTOIOl
;
else
assign
CAHBLTIIIOl
=
1
'b
0
;
if
(
CAHBLTlIO0
[
10
]
)
assign
CAHBLTlIIOl
=
CAHBLTOIOl
;
else
assign
CAHBLTlIIOl
=
1
'b
0
;
if
(
CAHBLTlIO0
[
11
]
)
assign
CAHBLTOlIOl
=
CAHBLTOIOl
;
else
assign
CAHBLTOlIOl
=
1
'b
0
;
if
(
CAHBLTlIO0
[
12
]
)
assign
CAHBLTIlIOl
=
CAHBLTOIOl
;
else
assign
CAHBLTIlIOl
=
1
'b
0
;
if
(
CAHBLTlIO0
[
13
]
)
assign
CAHBLTllIOl
=
CAHBLTOIOl
;
else
assign
CAHBLTllIOl
=
1
'b
0
;
if
(
CAHBLTlIO0
[
14
]
)
assign
CAHBLTO0IOl
=
CAHBLTOIOl
;
else
assign
CAHBLTO0IOl
=
1
'b
0
;
if
(
CAHBLTlIO0
[
15
]
)
assign
CAHBLTI0IOl
=
CAHBLTOIOl
;
else
assign
CAHBLTI0IOl
=
1
'b
0
;
if
(
CAHBLTlIO0
[
16
]
)
assign
CAHBLTl0IOl
=
CAHBLTOIOl
;
else
assign
CAHBLTl0IOl
=
1
'b
0
;
if
(
CAHBLTlIlll
[
0
]
)
assign
CAHBLTlI100
=
CAHBLTIlOl
;
else
assign
CAHBLTlI100
=
1
'b
0
;
if
(
CAHBLTlIlll
[
1
]
)
assign
CAHBLTOl100
=
CAHBLTIlOl
;
else
assign
CAHBLTOl100
=
1
'b
0
;
if
(
CAHBLTlIlll
[
2
]
)
assign
CAHBLTIl100
=
CAHBLTIlOl
;
else
assign
CAHBLTIl100
=
1
'b
0
;
if
(
CAHBLTlIlll
[
3
]
)
assign
CAHBLTll100
=
CAHBLTIlOl
;
else
assign
CAHBLTll100
=
1
'b
0
;
if
(
CAHBLTlIlll
[
4
]
)
assign
CAHBLTO0100
=
CAHBLTIlOl
;
else
assign
CAHBLTO0100
=
1
'b
0
;
if
(
CAHBLTlIlll
[
5
]
)
assign
CAHBLTI0100
=
CAHBLTIlOl
;
else
assign
CAHBLTI0100
=
1
'b
0
;
if
(
CAHBLTlIlll
[
6
]
)
assign
CAHBLTl0100
=
CAHBLTIlOl
;
else
assign
CAHBLTl0100
=
1
'b
0
;
if
(
CAHBLTlIlll
[
7
]
)
assign
CAHBLTO1100
=
CAHBLTIlOl
;
else
assign
CAHBLTO1100
=
1
'b
0
;
if
(
CAHBLTlIlll
[
8
]
)
assign
CAHBLTI1100
=
CAHBLTIlOl
;
else
assign
CAHBLTI1100
=
1
'b
0
;
if
(
CAHBLTlIlll
[
9
]
)
assign
CAHBLTl1100
=
CAHBLTIlOl
;
else
assign
CAHBLTl1100
=
1
'b
0
;
if
(
CAHBLTlIlll
[
10
]
)
assign
CAHBLTOOO10
=
CAHBLTIlOl
;
else
assign
CAHBLTOOO10
=
1
'b
0
;
if
(
CAHBLTlIlll
[
11
]
)
assign
CAHBLTIOO10
=
CAHBLTIlOl
;
else
assign
CAHBLTIOO10
=
1
'b
0
;
if
(
CAHBLTlIlll
[
12
]
)
assign
CAHBLTlOO10
=
CAHBLTIlOl
;
else
assign
CAHBLTlOO10
=
1
'b
0
;
if
(
CAHBLTlIlll
[
13
]
)
assign
CAHBLTOIO10
=
CAHBLTIlOl
;
else
assign
CAHBLTOIO10
=
1
'b
0
;
if
(
CAHBLTlIlll
[
14
]
)
assign
CAHBLTIIO10
=
CAHBLTIlOl
;
else
assign
CAHBLTIIO10
=
1
'b
0
;
if
(
CAHBLTlIlll
[
15
]
)
assign
CAHBLTlIO10
=
CAHBLTIlOl
;
else
assign
CAHBLTlIO10
=
1
'b
0
;
if
(
CAHBLTlIlll
[
16
]
)
assign
CAHBLTOlO10
=
CAHBLTIlOl
;
else
assign
CAHBLTOlO10
=
1
'b
0
;
if
(
CAHBLTOllll
[
0
]
)
assign
CAHBLTIlO10
=
CAHBLTl0Ol
;
else
assign
CAHBLTIlO10
=
1
'b
0
;
if
(
CAHBLTOllll
[
1
]
)
assign
CAHBLTllO10
=
CAHBLTl0Ol
;
else
assign
CAHBLTllO10
=
1
'b
0
;
if
(
CAHBLTOllll
[
2
]
)
assign
CAHBLTO0O10
=
CAHBLTl0Ol
;
else
assign
CAHBLTO0O10
=
1
'b
0
;
if
(
CAHBLTOllll
[
3
]
)
assign
CAHBLTI0O10
=
CAHBLTl0Ol
;
else
assign
CAHBLTI0O10
=
1
'b
0
;
if
(
CAHBLTOllll
[
4
]
)
assign
CAHBLTl0O10
=
CAHBLTl0Ol
;
else
assign
CAHBLTl0O10
=
1
'b
0
;
if
(
CAHBLTOllll
[
5
]
)
assign
CAHBLTO1O10
=
CAHBLTl0Ol
;
else
assign
CAHBLTO1O10
=
1
'b
0
;
if
(
CAHBLTOllll
[
6
]
)
assign
CAHBLTI1O10
=
CAHBLTl0Ol
;
else
assign
CAHBLTI1O10
=
1
'b
0
;
if
(
CAHBLTOllll
[
7
]
)
assign
CAHBLTl1O10
=
CAHBLTl0Ol
;
else
assign
CAHBLTl1O10
=
1
'b
0
;
if
(
CAHBLTOllll
[
8
]
)
assign
CAHBLTOOI10
=
CAHBLTl0Ol
;
else
assign
CAHBLTOOI10
=
1
'b
0
;
if
(
CAHBLTOllll
[
9
]
)
assign
CAHBLTIOI10
=
CAHBLTl0Ol
;
else
assign
CAHBLTIOI10
=
1
'b
0
;
if
(
CAHBLTOllll
[
10
]
)
assign
CAHBLTlOI10
=
CAHBLTl0Ol
;
else
assign
CAHBLTlOI10
=
1
'b
0
;
if
(
CAHBLTOllll
[
11
]
)
assign
CAHBLTOII10
=
CAHBLTl0Ol
;
else
assign
CAHBLTOII10
=
1
'b
0
;
if
(
CAHBLTOllll
[
12
]
)
assign
CAHBLTIII10
=
CAHBLTl0Ol
;
else
assign
CAHBLTIII10
=
1
'b
0
;
if
(
CAHBLTOllll
[
13
]
)
assign
CAHBLTlII10
=
CAHBLTl0Ol
;
else
assign
CAHBLTlII10
=
1
'b
0
;
if
(
CAHBLTOllll
[
14
]
)
assign
CAHBLTOlI10
=
CAHBLTl0Ol
;
else
assign
CAHBLTOlI10
=
1
'b
0
;
if
(
CAHBLTOllll
[
15
]
)
assign
CAHBLTIlI10
=
CAHBLTl0Ol
;
else
assign
CAHBLTIlI10
=
1
'b
0
;
if
(
CAHBLTOllll
[
16
]
)
assign
CAHBLTllI10
=
CAHBLTl0Ol
;
else
assign
CAHBLTllI10
=
1
'b
0
;
endgenerate
generate
if
(
CAHBLTIIO0
[
0
]
)
assign
CAHBLTIO1Ol
=
CAHBLTOOOl
;
else
assign
CAHBLTIO1Ol
=
1
'b
0
;
if
(
CAHBLTIIO0
[
1
]
)
assign
CAHBLTlO1Ol
=
CAHBLTOOOl
;
else
assign
CAHBLTlO1Ol
=
1
'b
0
;
if
(
CAHBLTIIO0
[
2
]
)
assign
CAHBLTOI1Ol
=
CAHBLTOOOl
;
else
assign
CAHBLTOI1Ol
=
1
'b
0
;
if
(
CAHBLTIIO0
[
3
]
)
assign
CAHBLTII1Ol
=
CAHBLTOOOl
;
else
assign
CAHBLTII1Ol
=
1
'b
0
;
if
(
CAHBLTIIO0
[
4
]
)
assign
CAHBLTlI1Ol
=
CAHBLTOOOl
;
else
assign
CAHBLTlI1Ol
=
1
'b
0
;
if
(
CAHBLTIIO0
[
5
]
)
assign
CAHBLTOl1Ol
=
CAHBLTOOOl
;
else
assign
CAHBLTOl1Ol
=
1
'b
0
;
if
(
CAHBLTIIO0
[
6
]
)
assign
CAHBLTIl1Ol
=
CAHBLTOOOl
;
else
assign
CAHBLTIl1Ol
=
1
'b
0
;
if
(
CAHBLTIIO0
[
7
]
)
assign
CAHBLTll1Ol
=
CAHBLTOOOl
;
else
assign
CAHBLTll1Ol
=
1
'b
0
;
if
(
CAHBLTIIO0
[
8
]
)
assign
CAHBLTO01Ol
=
CAHBLTOOOl
;
else
assign
CAHBLTO01Ol
=
1
'b
0
;
if
(
CAHBLTIIO0
[
9
]
)
assign
CAHBLTI01Ol
=
CAHBLTOOOl
;
else
assign
CAHBLTI01Ol
=
1
'b
0
;
if
(
CAHBLTIIO0
[
10
]
)
assign
CAHBLTl01Ol
=
CAHBLTOOOl
;
else
assign
CAHBLTl01Ol
=
1
'b
0
;
if
(
CAHBLTIIO0
[
11
]
)
assign
CAHBLTO11Ol
=
CAHBLTOOOl
;
else
assign
CAHBLTO11Ol
=
1
'b
0
;
if
(
CAHBLTIIO0
[
12
]
)
assign
CAHBLTI11Ol
=
CAHBLTOOOl
;
else
assign
CAHBLTI11Ol
=
1
'b
0
;
if
(
CAHBLTIIO0
[
13
]
)
assign
CAHBLTl11Ol
=
CAHBLTOOOl
;
else
assign
CAHBLTl11Ol
=
1
'b
0
;
if
(
CAHBLTIIO0
[
14
]
)
assign
CAHBLTOOOIl
=
CAHBLTOOOl
;
else
assign
CAHBLTOOOIl
=
1
'b
0
;
if
(
CAHBLTIIO0
[
15
]
)
assign
CAHBLTIOOIl
=
CAHBLTOOOl
;
else
assign
CAHBLTIOOIl
=
1
'b
0
;
if
(
CAHBLTIIO0
[
16
]
)
assign
CAHBLTlOOIl
=
CAHBLTOOOl
;
else
assign
CAHBLTlOOIl
=
1
'b
0
;
if
(
CAHBLTlIO0
[
0
]
)
assign
CAHBLTOIOIl
=
CAHBLTIIOl
;
else
assign
CAHBLTOIOIl
=
1
'b
0
;
if
(
CAHBLTlIO0
[
1
]
)
assign
CAHBLTIIOIl
=
CAHBLTIIOl
;
else
assign
CAHBLTIIOIl
=
1
'b
0
;
if
(
CAHBLTlIO0
[
2
]
)
assign
CAHBLTlIOIl
=
CAHBLTIIOl
;
else
assign
CAHBLTlIOIl
=
1
'b
0
;
if
(
CAHBLTlIO0
[
3
]
)
assign
CAHBLTOlOIl
=
CAHBLTIIOl
;
else
assign
CAHBLTOlOIl
=
1
'b
0
;
if
(
CAHBLTlIO0
[
4
]
)
assign
CAHBLTIlOIl
=
CAHBLTIIOl
;
else
assign
CAHBLTIlOIl
=
1
'b
0
;
if
(
CAHBLTlIO0
[
5
]
)
assign
CAHBLTllOIl
=
CAHBLTIIOl
;
else
assign
CAHBLTllOIl
=
1
'b
0
;
if
(
CAHBLTlIO0
[
6
]
)
assign
CAHBLTO0OIl
=
CAHBLTIIOl
;
else
assign
CAHBLTO0OIl
=
1
'b
0
;
if
(
CAHBLTlIO0
[
7
]
)
assign
CAHBLTI0OIl
=
CAHBLTIIOl
;
else
assign
CAHBLTI0OIl
=
1
'b
0
;
if
(
CAHBLTlIO0
[
8
]
)
assign
CAHBLTl0OIl
=
CAHBLTIIOl
;
else
assign
CAHBLTl0OIl
=
1
'b
0
;
if
(
CAHBLTlIO0
[
9
]
)
assign
CAHBLTO1OIl
=
CAHBLTIIOl
;
else
assign
CAHBLTO1OIl
=
1
'b
0
;
if
(
CAHBLTlIO0
[
10
]
)
assign
CAHBLTI1OIl
=
CAHBLTIIOl
;
else
assign
CAHBLTI1OIl
=
1
'b
0
;
if
(
CAHBLTlIO0
[
11
]
)
assign
CAHBLTl1OIl
=
CAHBLTIIOl
;
else
assign
CAHBLTl1OIl
=
1
'b
0
;
if
(
CAHBLTlIO0
[
12
]
)
assign
CAHBLTOOIIl
=
CAHBLTIIOl
;
else
assign
CAHBLTOOIIl
=
1
'b
0
;
if
(
CAHBLTlIO0
[
13
]
)
assign
CAHBLTIOIIl
=
CAHBLTIIOl
;
else
assign
CAHBLTIOIIl
=
1
'b
0
;
if
(
CAHBLTlIO0
[
14
]
)
assign
CAHBLTlOIIl
=
CAHBLTIIOl
;
else
assign
CAHBLTlOIIl
=
1
'b
0
;
if
(
CAHBLTlIO0
[
15
]
)
assign
CAHBLTOIIIl
=
CAHBLTIIOl
;
else
assign
CAHBLTOIIIl
=
1
'b
0
;
if
(
CAHBLTlIO0
[
16
]
)
assign
CAHBLTIIIIl
=
CAHBLTIIOl
;
else
assign
CAHBLTIIIIl
=
1
'b
0
;
if
(
CAHBLTlIlll
[
0
]
)
assign
CAHBLTI1010
=
CAHBLTllOl
;
else
assign
CAHBLTI1010
=
1
'b
0
;
if
(
CAHBLTlIlll
[
1
]
)
assign
CAHBLTl1010
=
CAHBLTllOl
;
else
assign
CAHBLTl1010
=
1
'b
0
;
if
(
CAHBLTlIlll
[
2
]
)
assign
CAHBLTOO110
=
CAHBLTllOl
;
else
assign
CAHBLTOO110
=
1
'b
0
;
if
(
CAHBLTlIlll
[
3
]
)
assign
CAHBLTIO110
=
CAHBLTllOl
;
else
assign
CAHBLTIO110
=
1
'b
0
;
if
(
CAHBLTlIlll
[
4
]
)
assign
CAHBLTlO110
=
CAHBLTllOl
;
else
assign
CAHBLTlO110
=
1
'b
0
;
if
(
CAHBLTlIlll
[
5
]
)
assign
CAHBLTOI110
=
CAHBLTllOl
;
else
assign
CAHBLTOI110
=
1
'b
0
;
if
(
CAHBLTlIlll
[
6
]
)
assign
CAHBLTII110
=
CAHBLTllOl
;
else
assign
CAHBLTII110
=
1
'b
0
;
if
(
CAHBLTlIlll
[
7
]
)
assign
CAHBLTlI110
=
CAHBLTllOl
;
else
assign
CAHBLTlI110
=
1
'b
0
;
if
(
CAHBLTlIlll
[
8
]
)
assign
CAHBLTOl110
=
CAHBLTllOl
;
else
assign
CAHBLTOl110
=
1
'b
0
;
if
(
CAHBLTlIlll
[
9
]
)
assign
CAHBLTIl110
=
CAHBLTllOl
;
else
assign
CAHBLTIl110
=
1
'b
0
;
if
(
CAHBLTlIlll
[
10
]
)
assign
CAHBLTll110
=
CAHBLTllOl
;
else
assign
CAHBLTll110
=
1
'b
0
;
if
(
CAHBLTlIlll
[
11
]
)
assign
CAHBLTO0110
=
CAHBLTllOl
;
else
assign
CAHBLTO0110
=
1
'b
0
;
if
(
CAHBLTlIlll
[
12
]
)
assign
CAHBLTI0110
=
CAHBLTllOl
;
else
assign
CAHBLTI0110
=
1
'b
0
;
if
(
CAHBLTlIlll
[
13
]
)
assign
CAHBLTl0110
=
CAHBLTllOl
;
else
assign
CAHBLTl0110
=
1
'b
0
;
if
(
CAHBLTlIlll
[
14
]
)
assign
CAHBLTO1110
=
CAHBLTllOl
;
else
assign
CAHBLTO1110
=
1
'b
0
;
if
(
CAHBLTlIlll
[
15
]
)
assign
CAHBLTI1110
=
CAHBLTllOl
;
else
assign
CAHBLTI1110
=
1
'b
0
;
if
(
CAHBLTlIlll
[
16
]
)
assign
CAHBLTl1110
=
CAHBLTllOl
;
else
assign
CAHBLTl1110
=
1
'b
0
;
if
(
CAHBLTOllll
[
0
]
)
assign
CAHBLTOOOO1
=
CAHBLTO1Ol
;
else
assign
CAHBLTOOOO1
=
1
'b
0
;
if
(
CAHBLTOllll
[
1
]
)
assign
CAHBLTIOOO1
=
CAHBLTO1Ol
;
else
assign
CAHBLTIOOO1
=
1
'b
0
;
if
(
CAHBLTOllll
[
2
]
)
assign
CAHBLTlOOO1
=
CAHBLTO1Ol
;
else
assign
CAHBLTlOOO1
=
1
'b
0
;
if
(
CAHBLTOllll
[
3
]
)
assign
CAHBLTOIOO1
=
CAHBLTO1Ol
;
else
assign
CAHBLTOIOO1
=
1
'b
0
;
if
(
CAHBLTOllll
[
4
]
)
assign
CAHBLTIIOO1
=
CAHBLTO1Ol
;
else
assign
CAHBLTIIOO1
=
1
'b
0
;
if
(
CAHBLTOllll
[
5
]
)
assign
CAHBLTlIOO1
=
CAHBLTO1Ol
;
else
assign
CAHBLTlIOO1
=
1
'b
0
;
if
(
CAHBLTOllll
[
6
]
)
assign
CAHBLTOlOO1
=
CAHBLTO1Ol
;
else
assign
CAHBLTOlOO1
=
1
'b
0
;
if
(
CAHBLTOllll
[
7
]
)
assign
CAHBLTIlOO1
=
CAHBLTO1Ol
;
else
assign
CAHBLTIlOO1
=
1
'b
0
;
if
(
CAHBLTOllll
[
8
]
)
assign
CAHBLTllOO1
=
CAHBLTO1Ol
;
else
assign
CAHBLTllOO1
=
1
'b
0
;
if
(
CAHBLTOllll
[
9
]
)
assign
CAHBLTO0OO1
=
CAHBLTO1Ol
;
else
assign
CAHBLTO0OO1
=
1
'b
0
;
if
(
CAHBLTOllll
[
10
]
)
assign
CAHBLTI0OO1
=
CAHBLTO1Ol
;
else
assign
CAHBLTI0OO1
=
1
'b
0
;
if
(
CAHBLTOllll
[
11
]
)
assign
CAHBLTl0OO1
=
CAHBLTO1Ol
;
else
assign
CAHBLTl0OO1
=
1
'b
0
;
if
(
CAHBLTOllll
[
12
]
)
assign
CAHBLTO1OO1
=
CAHBLTO1Ol
;
else
assign
CAHBLTO1OO1
=
1
'b
0
;
if
(
CAHBLTOllll
[
13
]
)
assign
CAHBLTI1OO1
=
CAHBLTO1Ol
;
else
assign
CAHBLTI1OO1
=
1
'b
0
;
if
(
CAHBLTOllll
[
14
]
)
assign
CAHBLTl1OO1
=
CAHBLTO1Ol
;
else
assign
CAHBLTl1OO1
=
1
'b
0
;
if
(
CAHBLTOllll
[
15
]
)
assign
CAHBLTOOIO1
=
CAHBLTO1Ol
;
else
assign
CAHBLTOOIO1
=
1
'b
0
;
if
(
CAHBLTOllll
[
16
]
)
assign
CAHBLTIOIO1
=
CAHBLTO1Ol
;
else
assign
CAHBLTIOIO1
=
1
'b
0
;
endgenerate
generate
if
(
CAHBLTIIO0
[
0
]
)
assign
CAHBLTlIIIl
=
CAHBLTIOOl
;
else
assign
CAHBLTlIIIl
=
1
'b
0
;
if
(
CAHBLTIIO0
[
1
]
)
assign
CAHBLTOlIIl
=
CAHBLTIOOl
;
else
assign
CAHBLTOlIIl
=
1
'b
0
;
if
(
CAHBLTIIO0
[
2
]
)
assign
CAHBLTIlIIl
=
CAHBLTIOOl
;
else
assign
CAHBLTIlIIl
=
1
'b
0
;
if
(
CAHBLTIIO0
[
3
]
)
assign
CAHBLTllIIl
=
CAHBLTIOOl
;
else
assign
CAHBLTllIIl
=
1
'b
0
;
if
(
CAHBLTIIO0
[
4
]
)
assign
CAHBLTO0IIl
=
CAHBLTIOOl
;
else
assign
CAHBLTO0IIl
=
1
'b
0
;
if
(
CAHBLTIIO0
[
5
]
)
assign
CAHBLTI0IIl
=
CAHBLTIOOl
;
else
assign
CAHBLTI0IIl
=
1
'b
0
;
if
(
CAHBLTIIO0
[
6
]
)
assign
CAHBLTl0IIl
=
CAHBLTIOOl
;
else
assign
CAHBLTl0IIl
=
1
'b
0
;
if
(
CAHBLTIIO0
[
7
]
)
assign
CAHBLTO1IIl
=
CAHBLTIOOl
;
else
assign
CAHBLTO1IIl
=
1
'b
0
;
if
(
CAHBLTIIO0
[
8
]
)
assign
CAHBLTI1IIl
=
CAHBLTIOOl
;
else
assign
CAHBLTI1IIl
=
1
'b
0
;
if
(
CAHBLTIIO0
[
9
]
)
assign
CAHBLTl1IIl
=
CAHBLTIOOl
;
else
assign
CAHBLTl1IIl
=
1
'b
0
;
if
(
CAHBLTIIO0
[
10
]
)
assign
CAHBLTOOlIl
=
CAHBLTIOOl
;
else
assign
CAHBLTOOlIl
=
1
'b
0
;
if
(
CAHBLTIIO0
[
11
]
)
assign
CAHBLTIOlIl
=
CAHBLTIOOl
;
else
assign
CAHBLTIOlIl
=
1
'b
0
;
if
(
CAHBLTIIO0
[
12
]
)
assign
CAHBLTlOlIl
=
CAHBLTIOOl
;
else
assign
CAHBLTlOlIl
=
1
'b
0
;
if
(
CAHBLTIIO0
[
13
]
)
assign
CAHBLTOIlIl
=
CAHBLTIOOl
;
else
assign
CAHBLTOIlIl
=
1
'b
0
;
if
(
CAHBLTIIO0
[
14
]
)
assign
CAHBLTIIlIl
=
CAHBLTIOOl
;
else
assign
CAHBLTIIlIl
=
1
'b
0
;
if
(
CAHBLTIIO0
[
15
]
)
assign
CAHBLTlIlIl
=
CAHBLTIOOl
;
else
assign
CAHBLTlIlIl
=
1
'b
0
;
if
(
CAHBLTIIO0
[
16
]
)
assign
CAHBLTOllIl
=
CAHBLTIOOl
;
else
assign
CAHBLTOllIl
=
1
'b
0
;
if
(
CAHBLTlIO0
[
0
]
)
assign
CAHBLTIllIl
=
CAHBLTlIOl
;
else
assign
CAHBLTIllIl
=
1
'b
0
;
if
(
CAHBLTlIO0
[
1
]
)
assign
CAHBLTlllIl
=
CAHBLTlIOl
;
else
assign
CAHBLTlllIl
=
1
'b
0
;
if
(
CAHBLTlIO0
[
2
]
)
assign
CAHBLTO0lIl
=
CAHBLTlIOl
;
else
assign
CAHBLTO0lIl
=
1
'b
0
;
if
(
CAHBLTlIO0
[
3
]
)
assign
CAHBLTI0lIl
=
CAHBLTlIOl
;
else
assign
CAHBLTI0lIl
=
1
'b
0
;
if
(
CAHBLTlIO0
[
4
]
)
assign
CAHBLTl0lIl
=
CAHBLTlIOl
;
else
assign
CAHBLTl0lIl
=
1
'b
0
;
if
(
CAHBLTlIO0
[
5
]
)
assign
CAHBLTO1lIl
=
CAHBLTlIOl
;
else
assign
CAHBLTO1lIl
=
1
'b
0
;
if
(
CAHBLTlIO0
[
6
]
)
assign
CAHBLTI1lIl
=
CAHBLTlIOl
;
else
assign
CAHBLTI1lIl
=
1
'b
0
;
if
(
CAHBLTlIO0
[
7
]
)
assign
CAHBLTl1lIl
=
CAHBLTlIOl
;
else
assign
CAHBLTl1lIl
=
1
'b
0
;
if
(
CAHBLTlIO0
[
8
]
)
assign
CAHBLTOO0Il
=
CAHBLTlIOl
;
else
assign
CAHBLTOO0Il
=
1
'b
0
;
if
(
CAHBLTlIO0
[
9
]
)
assign
CAHBLTIO0Il
=
CAHBLTlIOl
;
else
assign
CAHBLTIO0Il
=
1
'b
0
;
if
(
CAHBLTlIO0
[
10
]
)
assign
CAHBLTlO0Il
=
CAHBLTlIOl
;
else
assign
CAHBLTlO0Il
=
1
'b
0
;
if
(
CAHBLTlIO0
[
11
]
)
assign
CAHBLTOI0Il
=
CAHBLTlIOl
;
else
assign
CAHBLTOI0Il
=
1
'b
0
;
if
(
CAHBLTlIO0
[
12
]
)
assign
CAHBLTII0Il
=
CAHBLTlIOl
;
else
assign
CAHBLTII0Il
=
1
'b
0
;
if
(
CAHBLTlIO0
[
13
]
)
assign
CAHBLTlI0Il
=
CAHBLTlIOl
;
else
assign
CAHBLTlI0Il
=
1
'b
0
;
if
(
CAHBLTlIO0
[
14
]
)
assign
CAHBLTOl0Il
=
CAHBLTlIOl
;
else
assign
CAHBLTOl0Il
=
1
'b
0
;
if
(
CAHBLTlIO0
[
15
]
)
assign
CAHBLTIl0Il
=
CAHBLTlIOl
;
else
assign
CAHBLTIl0Il
=
1
'b
0
;
if
(
CAHBLTlIO0
[
16
]
)
assign
CAHBLTll0Il
=
CAHBLTlIOl
;
else
assign
CAHBLTll0Il
=
1
'b
0
;
if
(
CAHBLTlIlll
[
0
]
)
assign
CAHBLTlOIO1
=
CAHBLTO0Ol
;
else
assign
CAHBLTlOIO1
=
1
'b
0
;
if
(
CAHBLTlIlll
[
1
]
)
assign
CAHBLTOIIO1
=
CAHBLTO0Ol
;
else
assign
CAHBLTOIIO1
=
1
'b
0
;
if
(
CAHBLTlIlll
[
2
]
)
assign
CAHBLTIIIO1
=
CAHBLTO0Ol
;
else
assign
CAHBLTIIIO1
=
1
'b
0
;
if
(
CAHBLTlIlll
[
3
]
)
assign
CAHBLTlIIO1
=
CAHBLTO0Ol
;
else
assign
CAHBLTlIIO1
=
1
'b
0
;
if
(
CAHBLTlIlll
[
4
]
)
assign
CAHBLTOlIO1
=
CAHBLTO0Ol
;
else
assign
CAHBLTOlIO1
=
1
'b
0
;
if
(
CAHBLTlIlll
[
5
]
)
assign
CAHBLTIlIO1
=
CAHBLTO0Ol
;
else
assign
CAHBLTIlIO1
=
1
'b
0
;
if
(
CAHBLTlIlll
[
6
]
)
assign
CAHBLTllIO1
=
CAHBLTO0Ol
;
else
assign
CAHBLTllIO1
=
1
'b
0
;
if
(
CAHBLTlIlll
[
7
]
)
assign
CAHBLTO0IO1
=
CAHBLTO0Ol
;
else
assign
CAHBLTO0IO1
=
1
'b
0
;
if
(
CAHBLTlIlll
[
8
]
)
assign
CAHBLTI0IO1
=
CAHBLTO0Ol
;
else
assign
CAHBLTI0IO1
=
1
'b
0
;
if
(
CAHBLTlIlll
[
9
]
)
assign
CAHBLTl0IO1
=
CAHBLTO0Ol
;
else
assign
CAHBLTl0IO1
=
1
'b
0
;
if
(
CAHBLTlIlll
[
10
]
)
assign
CAHBLTO1IO1
=
CAHBLTO0Ol
;
else
assign
CAHBLTO1IO1
=
1
'b
0
;
if
(
CAHBLTlIlll
[
11
]
)
assign
CAHBLTI1IO1
=
CAHBLTO0Ol
;
else
assign
CAHBLTI1IO1
=
1
'b
0
;
if
(
CAHBLTlIlll
[
12
]
)
assign
CAHBLTl1IO1
=
CAHBLTO0Ol
;
else
assign
CAHBLTl1IO1
=
1
'b
0
;
if
(
CAHBLTlIlll
[
13
]
)
assign
CAHBLTOOlO1
=
CAHBLTO0Ol
;
else
assign
CAHBLTOOlO1
=
1
'b
0
;
if
(
CAHBLTlIlll
[
14
]
)
assign
CAHBLTIOlO1
=
CAHBLTO0Ol
;
else
assign
CAHBLTIOlO1
=
1
'b
0
;
if
(
CAHBLTlIlll
[
15
]
)
assign
CAHBLTlOlO1
=
CAHBLTO0Ol
;
else
assign
CAHBLTlOlO1
=
1
'b
0
;
if
(
CAHBLTlIlll
[
16
]
)
assign
CAHBLTOIlO1
=
CAHBLTO0Ol
;
else
assign
CAHBLTOIlO1
=
1
'b
0
;
if
(
CAHBLTOllll
[
0
]
)
assign
CAHBLTIIlO1
=
CAHBLTI1Ol
;
else
assign
CAHBLTIIlO1
=
1
'b
0
;
if
(
CAHBLTOllll
[
1
]
)
assign
CAHBLTlIlO1
=
CAHBLTI1Ol
;
else
assign
CAHBLTlIlO1
=
1
'b
0
;
if
(
CAHBLTOllll
[
2
]
)
assign
CAHBLTOllO1
=
CAHBLTI1Ol
;
else
assign
CAHBLTOllO1
=
1
'b
0
;
if
(
CAHBLTOllll
[
3
]
)
assign
CAHBLTIllO1
=
CAHBLTI1Ol
;
else
assign
CAHBLTIllO1
=
1
'b
0
;
if
(
CAHBLTOllll
[
4
]
)
assign
CAHBLTlllO1
=
CAHBLTI1Ol
;
else
assign
CAHBLTlllO1
=
1
'b
0
;
if
(
CAHBLTOllll
[
5
]
)
assign
CAHBLTO0lO1
=
CAHBLTI1Ol
;
else
assign
CAHBLTO0lO1
=
1
'b
0
;
if
(
CAHBLTOllll
[
6
]
)
assign
CAHBLTI0lO1
=
CAHBLTI1Ol
;
else
assign
CAHBLTI0lO1
=
1
'b
0
;
if
(
CAHBLTOllll
[
7
]
)
assign
CAHBLTl0lO1
=
CAHBLTI1Ol
;
else
assign
CAHBLTl0lO1
=
1
'b
0
;
if
(
CAHBLTOllll
[
8
]
)
assign
CAHBLTO1lO1
=
CAHBLTI1Ol
;
else
assign
CAHBLTO1lO1
=
1
'b
0
;
if
(
CAHBLTOllll
[
9
]
)
assign
CAHBLTI1lO1
=
CAHBLTI1Ol
;
else
assign
CAHBLTI1lO1
=
1
'b
0
;
if
(
CAHBLTOllll
[
10
]
)
assign
CAHBLTl1lO1
=
CAHBLTI1Ol
;
else
assign
CAHBLTl1lO1
=
1
'b
0
;
if
(
CAHBLTOllll
[
11
]
)
assign
CAHBLTOO0O1
=
CAHBLTI1Ol
;
else
assign
CAHBLTOO0O1
=
1
'b
0
;
if
(
CAHBLTOllll
[
12
]
)
assign
CAHBLTIO0O1
=
CAHBLTI1Ol
;
else
assign
CAHBLTIO0O1
=
1
'b
0
;
if
(
CAHBLTOllll
[
13
]
)
assign
CAHBLTlO0O1
=
CAHBLTI1Ol
;
else
assign
CAHBLTlO0O1
=
1
'b
0
;
if
(
CAHBLTOllll
[
14
]
)
assign
CAHBLTOI0O1
=
CAHBLTI1Ol
;
else
assign
CAHBLTOI0O1
=
1
'b
0
;
if
(
CAHBLTOllll
[
15
]
)
assign
CAHBLTII0O1
=
CAHBLTI1Ol
;
else
assign
CAHBLTII0O1
=
1
'b
0
;
if
(
CAHBLTOllll
[
16
]
)
assign
CAHBLTlI0O1
=
CAHBLTI1Ol
;
else
assign
CAHBLTlI0O1
=
1
'b
0
;
endgenerate
generate
if
(
CAHBLTIIO0
[
0
]
)
assign
CAHBLTO00Il
=
CAHBLTOlO0
;
else
assign
CAHBLTO00Il
=
1
'b
1
;
if
(
CAHBLTIIO0
[
1
]
)
assign
CAHBLTI00Il
=
CAHBLTOlO0
;
else
assign
CAHBLTI00Il
=
1
'b
1
;
if
(
CAHBLTIIO0
[
2
]
)
assign
CAHBLTl00Il
=
CAHBLTOlO0
;
else
assign
CAHBLTl00Il
=
1
'b
1
;
if
(
CAHBLTIIO0
[
3
]
)
assign
CAHBLTO10Il
=
CAHBLTOlO0
;
else
assign
CAHBLTO10Il
=
1
'b
1
;
if
(
CAHBLTIIO0
[
4
]
)
assign
CAHBLTI10Il
=
CAHBLTOlO0
;
else
assign
CAHBLTI10Il
=
1
'b
1
;
if
(
CAHBLTIIO0
[
5
]
)
assign
CAHBLTl10Il
=
CAHBLTOlO0
;
else
assign
CAHBLTl10Il
=
1
'b
1
;
if
(
CAHBLTIIO0
[
6
]
)
assign
CAHBLTOO1Il
=
CAHBLTOlO0
;
else
assign
CAHBLTOO1Il
=
1
'b
1
;
if
(
CAHBLTIIO0
[
7
]
)
assign
CAHBLTIO1Il
=
CAHBLTOlO0
;
else
assign
CAHBLTIO1Il
=
1
'b
1
;
if
(
CAHBLTIIO0
[
8
]
)
assign
CAHBLTlO1Il
=
CAHBLTOlO0
;
else
assign
CAHBLTlO1Il
=
1
'b
1
;
if
(
CAHBLTIIO0
[
9
]
)
assign
CAHBLTOI1Il
=
CAHBLTOlO0
;
else
assign
CAHBLTOI1Il
=
1
'b
1
;
if
(
CAHBLTIIO0
[
10
]
)
assign
CAHBLTII1Il
=
CAHBLTOlO0
;
else
assign
CAHBLTII1Il
=
1
'b
1
;
if
(
CAHBLTIIO0
[
11
]
)
assign
CAHBLTlI1Il
=
CAHBLTOlO0
;
else
assign
CAHBLTlI1Il
=
1
'b
1
;
if
(
CAHBLTIIO0
[
12
]
)
assign
CAHBLTOl1Il
=
CAHBLTOlO0
;
else
assign
CAHBLTOl1Il
=
1
'b
1
;
if
(
CAHBLTIIO0
[
13
]
)
assign
CAHBLTIl1Il
=
CAHBLTOlO0
;
else
assign
CAHBLTIl1Il
=
1
'b
1
;
if
(
CAHBLTIIO0
[
14
]
)
assign
CAHBLTll1Il
=
CAHBLTOlO0
;
else
assign
CAHBLTll1Il
=
1
'b
1
;
if
(
CAHBLTIIO0
[
15
]
)
assign
CAHBLTO01Il
=
CAHBLTOlO0
;
else
assign
CAHBLTO01Il
=
1
'b
1
;
if
(
CAHBLTIIO0
[
16
]
)
assign
CAHBLTI01Il
=
CAHBLTOlO0
;
else
assign
CAHBLTI01Il
=
1
'b
1
;
if
(
CAHBLTlIO0
[
0
]
)
assign
CAHBLTl01Il
=
CAHBLTO1IOI
;
else
assign
CAHBLTl01Il
=
1
'b
1
;
if
(
CAHBLTlIO0
[
1
]
)
assign
CAHBLTO11Il
=
CAHBLTO1IOI
;
else
assign
CAHBLTO11Il
=
1
'b
1
;
if
(
CAHBLTlIO0
[
2
]
)
assign
CAHBLTI11Il
=
CAHBLTO1IOI
;
else
assign
CAHBLTI11Il
=
1
'b
1
;
if
(
CAHBLTlIO0
[
3
]
)
assign
CAHBLTl11Il
=
CAHBLTO1IOI
;
else
assign
CAHBLTl11Il
=
1
'b
1
;
if
(
CAHBLTlIO0
[
4
]
)
assign
CAHBLTOOOll
=
CAHBLTO1IOI
;
else
assign
CAHBLTOOOll
=
1
'b
1
;
if
(
CAHBLTlIO0
[
5
]
)
assign
CAHBLTIOOll
=
CAHBLTO1IOI
;
else
assign
CAHBLTIOOll
=
1
'b
1
;
if
(
CAHBLTlIO0
[
6
]
)
assign
CAHBLTlOOll
=
CAHBLTO1IOI
;
else
assign
CAHBLTlOOll
=
1
'b
1
;
if
(
CAHBLTlIO0
[
7
]
)
assign
CAHBLTOIOll
=
CAHBLTO1IOI
;
else
assign
CAHBLTOIOll
=
1
'b
1
;
if
(
CAHBLTlIO0
[
8
]
)
assign
CAHBLTIIOll
=
CAHBLTO1IOI
;
else
assign
CAHBLTIIOll
=
1
'b
1
;
if
(
CAHBLTlIO0
[
9
]
)
assign
CAHBLTlIOll
=
CAHBLTO1IOI
;
else
assign
CAHBLTlIOll
=
1
'b
1
;
if
(
CAHBLTlIO0
[
10
]
)
assign
CAHBLTOlOll
=
CAHBLTO1IOI
;
else
assign
CAHBLTOlOll
=
1
'b
1
;
if
(
CAHBLTlIO0
[
11
]
)
assign
CAHBLTIlOll
=
CAHBLTO1IOI
;
else
assign
CAHBLTIlOll
=
1
'b
1
;
if
(
CAHBLTlIO0
[
12
]
)
assign
CAHBLTllOll
=
CAHBLTO1IOI
;
else
assign
CAHBLTllOll
=
1
'b
1
;
if
(
CAHBLTlIO0
[
13
]
)
assign
CAHBLTO0Oll
=
CAHBLTO1IOI
;
else
assign
CAHBLTO0Oll
=
1
'b
1
;
if
(
CAHBLTlIO0
[
14
]
)
assign
CAHBLTI0Oll
=
CAHBLTO1IOI
;
else
assign
CAHBLTI0Oll
=
1
'b
1
;
if
(
CAHBLTlIO0
[
15
]
)
assign
CAHBLTl0Oll
=
CAHBLTO1IOI
;
else
assign
CAHBLTl0Oll
=
1
'b
1
;
if
(
CAHBLTlIO0
[
16
]
)
assign
CAHBLTO1Oll
=
CAHBLTO1IOI
;
else
assign
CAHBLTO1Oll
=
1
'b
1
;
if
(
CAHBLTlIlll
[
0
]
)
assign
CAHBLTOl0O1
=
CAHBLTIllll
;
else
assign
CAHBLTOl0O1
=
1
'b
1
;
if
(
CAHBLTlIlll
[
1
]
)
assign
CAHBLTIl0O1
=
CAHBLTIllll
;
else
assign
CAHBLTIl0O1
=
1
'b
1
;
if
(
CAHBLTlIlll
[
2
]
)
assign
CAHBLTll0O1
=
CAHBLTIllll
;
else
assign
CAHBLTll0O1
=
1
'b
1
;
if
(
CAHBLTlIlll
[
3
]
)
assign
CAHBLTO00O1
=
CAHBLTIllll
;
else
assign
CAHBLTO00O1
=
1
'b
1
;
if
(
CAHBLTlIlll
[
4
]
)
assign
CAHBLTI00O1
=
CAHBLTIllll
;
else
assign
CAHBLTI00O1
=
1
'b
1
;
if
(
CAHBLTlIlll
[
5
]
)
assign
CAHBLTl00O1
=
CAHBLTIllll
;
else
assign
CAHBLTl00O1
=
1
'b
1
;
if
(
CAHBLTlIlll
[
6
]
)
assign
CAHBLTO10O1
=
CAHBLTIllll
;
else
assign
CAHBLTO10O1
=
1
'b
1
;
if
(
CAHBLTlIlll
[
7
]
)
assign
CAHBLTI10O1
=
CAHBLTIllll
;
else
assign
CAHBLTI10O1
=
1
'b
1
;
if
(
CAHBLTlIlll
[
8
]
)
assign
CAHBLTl10O1
=
CAHBLTIllll
;
else
assign
CAHBLTl10O1
=
1
'b
1
;
if
(
CAHBLTlIlll
[
9
]
)
assign
CAHBLTOO1O1
=
CAHBLTIllll
;
else
assign
CAHBLTOO1O1
=
1
'b
1
;
if
(
CAHBLTlIlll
[
10
]
)
assign
CAHBLTIO1O1
=
CAHBLTIllll
;
else
assign
CAHBLTIO1O1
=
1
'b
1
;
if
(
CAHBLTlIlll
[
11
]
)
assign
CAHBLTlO1O1
=
CAHBLTIllll
;
else
assign
CAHBLTlO1O1
=
1
'b
1
;
if
(
CAHBLTlIlll
[
12
]
)
assign
CAHBLTOI1O1
=
CAHBLTIllll
;
else
assign
CAHBLTOI1O1
=
1
'b
1
;
if
(
CAHBLTlIlll
[
13
]
)
assign
CAHBLTII1O1
=
CAHBLTIllll
;
else
assign
CAHBLTII1O1
=
1
'b
1
;
if
(
CAHBLTlIlll
[
14
]
)
assign
CAHBLTlI1O1
=
CAHBLTIllll
;
else
assign
CAHBLTlI1O1
=
1
'b
1
;
if
(
CAHBLTlIlll
[
15
]
)
assign
CAHBLTOl1O1
=
CAHBLTIllll
;
else
assign
CAHBLTOl1O1
=
1
'b
1
;
if
(
CAHBLTlIlll
[
16
]
)
assign
CAHBLTIl1O1
=
CAHBLTIllll
;
else
assign
CAHBLTIl1O1
=
1
'b
1
;
if
(
CAHBLTOllll
[
0
]
)
assign
CAHBLTll1O1
=
CAHBLTI101l
;
else
assign
CAHBLTll1O1
=
1
'b
1
;
if
(
CAHBLTOllll
[
1
]
)
assign
CAHBLTO01O1
=
CAHBLTI101l
;
else
assign
CAHBLTO01O1
=
1
'b
1
;
if
(
CAHBLTOllll
[
2
]
)
assign
CAHBLTI01O1
=
CAHBLTI101l
;
else
assign
CAHBLTI01O1
=
1
'b
1
;
if
(
CAHBLTOllll
[
3
]
)
assign
CAHBLTl01O1
=
CAHBLTI101l
;
else
assign
CAHBLTl01O1
=
1
'b
1
;
if
(
CAHBLTOllll
[
4
]
)
assign
CAHBLTO11O1
=
CAHBLTI101l
;
else
assign
CAHBLTO11O1
=
1
'b
1
;
if
(
CAHBLTOllll
[
5
]
)
assign
CAHBLTI11O1
=
CAHBLTI101l
;
else
assign
CAHBLTI11O1
=
1
'b
1
;
if
(
CAHBLTOllll
[
6
]
)
assign
CAHBLTl11O1
=
CAHBLTI101l
;
else
assign
CAHBLTl11O1
=
1
'b
1
;
if
(
CAHBLTOllll
[
7
]
)
assign
CAHBLTOOOI1
=
CAHBLTI101l
;
else
assign
CAHBLTOOOI1
=
1
'b
1
;
if
(
CAHBLTOllll
[
8
]
)
assign
CAHBLTIOOI1
=
CAHBLTI101l
;
else
assign
CAHBLTIOOI1
=
1
'b
1
;
if
(
CAHBLTOllll
[
9
]
)
assign
CAHBLTlOOI1
=
CAHBLTI101l
;
else
assign
CAHBLTlOOI1
=
1
'b
1
;
if
(
CAHBLTOllll
[
10
]
)
assign
CAHBLTOIOI1
=
CAHBLTI101l
;
else
assign
CAHBLTOIOI1
=
1
'b
1
;
if
(
CAHBLTOllll
[
11
]
)
assign
CAHBLTIIOI1
=
CAHBLTI101l
;
else
assign
CAHBLTIIOI1
=
1
'b
1
;
if
(
CAHBLTOllll
[
12
]
)
assign
CAHBLTlIOI1
=
CAHBLTI101l
;
else
assign
CAHBLTlIOI1
=
1
'b
1
;
if
(
CAHBLTOllll
[
13
]
)
assign
CAHBLTOlOI1
=
CAHBLTI101l
;
else
assign
CAHBLTOlOI1
=
1
'b
1
;
if
(
CAHBLTOllll
[
14
]
)
assign
CAHBLTIlOI1
=
CAHBLTI101l
;
else
assign
CAHBLTIlOI1
=
1
'b
1
;
if
(
CAHBLTOllll
[
15
]
)
assign
CAHBLTllOI1
=
CAHBLTI101l
;
else
assign
CAHBLTllOI1
=
1
'b
1
;
if
(
CAHBLTOllll
[
16
]
)
assign
CAHBLTO0OI1
=
CAHBLTI101l
;
else
assign
CAHBLTO0OI1
=
1
'b
1
;
endgenerate
generate
if
(
CAHBLTIIO0
[
0
]
)
assign
CAHBLTOI0lI
=
HRDATA_S0
;
else
assign
CAHBLTOI0lI
=
32
'h
0
;
if
(
CAHBLTIIO0
[
1
]
)
assign
CAHBLTII0lI
=
HRDATA_S1
;
else
assign
CAHBLTII0lI
=
32
'h
0
;
if
(
CAHBLTIIO0
[
2
]
)
assign
CAHBLTlI0lI
=
HRDATA_S2
;
else
assign
CAHBLTlI0lI
=
32
'h
0
;
if
(
CAHBLTIIO0
[
3
]
)
assign
CAHBLTOl0lI
=
HRDATA_S3
;
else
assign
CAHBLTOl0lI
=
32
'h
0
;
if
(
CAHBLTIIO0
[
4
]
)
assign
CAHBLTIl0lI
=
HRDATA_S4
;
else
assign
CAHBLTIl0lI
=
32
'h
0
;
if
(
CAHBLTIIO0
[
5
]
)
assign
CAHBLTll0lI
=
HRDATA_S5
;
else
assign
CAHBLTll0lI
=
32
'h
0
;
if
(
CAHBLTIIO0
[
6
]
)
assign
CAHBLTO00lI
=
HRDATA_S6
;
else
assign
CAHBLTO00lI
=
32
'h
0
;
if
(
CAHBLTIIO0
[
7
]
)
assign
CAHBLTI00lI
=
HRDATA_S7
;
else
assign
CAHBLTI00lI
=
32
'h
0
;
if
(
CAHBLTIIO0
[
8
]
)
assign
CAHBLTl00lI
=
HRDATA_S8
;
else
assign
CAHBLTl00lI
=
32
'h
0
;
if
(
CAHBLTIIO0
[
9
]
)
assign
CAHBLTO10lI
=
HRDATA_S9
;
else
assign
CAHBLTO10lI
=
32
'h
0
;
if
(
CAHBLTIIO0
[
10
]
)
assign
CAHBLTI10lI
=
HRDATA_S10
;
else
assign
CAHBLTI10lI
=
32
'h
0
;
if
(
CAHBLTIIO0
[
11
]
)
assign
CAHBLTl10lI
=
HRDATA_S11
;
else
assign
CAHBLTl10lI
=
32
'h
0
;
if
(
CAHBLTIIO0
[
12
]
)
assign
CAHBLTOO1lI
=
HRDATA_S12
;
else
assign
CAHBLTOO1lI
=
32
'h
0
;
if
(
CAHBLTIIO0
[
13
]
)
assign
CAHBLTIO1lI
=
HRDATA_S13
;
else
assign
CAHBLTIO1lI
=
32
'h
0
;
if
(
CAHBLTIIO0
[
14
]
)
assign
CAHBLTlO1lI
=
HRDATA_S14
;
else
assign
CAHBLTlO1lI
=
32
'h
0
;
if
(
CAHBLTIIO0
[
15
]
)
assign
CAHBLTOI1lI
=
HRDATA_S15
;
else
assign
CAHBLTOI1lI
=
32
'h
0
;
if
(
CAHBLTIIO0
[
16
]
)
assign
CAHBLTII1lI
=
HRDATA_S16
;
else
assign
CAHBLTII1lI
=
32
'h
0
;
if
(
CAHBLTlIO0
[
0
]
)
assign
CAHBLTlI1lI
=
HRDATA_S0
;
else
assign
CAHBLTlI1lI
=
32
'h
0
;
if
(
CAHBLTlIO0
[
1
]
)
assign
CAHBLTOl1lI
=
HRDATA_S1
;
else
assign
CAHBLTOl1lI
=
32
'h
0
;
if
(
CAHBLTlIO0
[
2
]
)
assign
CAHBLTIl1lI
=
HRDATA_S2
;
else
assign
CAHBLTIl1lI
=
32
'h
0
;
if
(
CAHBLTlIO0
[
3
]
)
assign
CAHBLTll1lI
=
HRDATA_S3
;
else
assign
CAHBLTll1lI
=
32
'h
0
;
if
(
CAHBLTlIO0
[
4
]
)
assign
CAHBLTO01lI
=
HRDATA_S4
;
else
assign
CAHBLTO01lI
=
32
'h
0
;
if
(
CAHBLTlIO0
[
5
]
)
assign
CAHBLTI01lI
=
HRDATA_S5
;
else
assign
CAHBLTI01lI
=
32
'h
0
;
if
(
CAHBLTlIO0
[
6
]
)
assign
CAHBLTl01lI
=
HRDATA_S6
;
else
assign
CAHBLTl01lI
=
32
'h
0
;
if
(
CAHBLTlIO0
[
7
]
)
assign
CAHBLTO11lI
=
HRDATA_S7
;
else
assign
CAHBLTO11lI
=
32
'h
0
;
if
(
CAHBLTlIO0
[
8
]
)
assign
CAHBLTI11lI
=
HRDATA_S8
;
else
assign
CAHBLTI11lI
=
32
'h
0
;
if
(
CAHBLTlIO0
[
9
]
)
assign
CAHBLTl11lI
=
HRDATA_S9
;
else
assign
CAHBLTl11lI
=
32
'h
0
;
if
(
CAHBLTlIO0
[
10
]
)
assign
CAHBLTOOO0I
=
HRDATA_S10
;
else
assign
CAHBLTOOO0I
=
32
'h
0
;
if
(
CAHBLTlIO0
[
11
]
)
assign
CAHBLTIOO0I
=
HRDATA_S11
;
else
assign
CAHBLTIOO0I
=
32
'h
0
;
if
(
CAHBLTlIO0
[
12
]
)
assign
CAHBLTlOO0I
=
HRDATA_S12
;
else
assign
CAHBLTlOO0I
=
32
'h
0
;
if
(
CAHBLTlIO0
[
13
]
)
assign
CAHBLTOIO0I
=
HRDATA_S13
;
else
assign
CAHBLTOIO0I
=
32
'h
0
;
if
(
CAHBLTlIO0
[
14
]
)
assign
CAHBLTIIO0I
=
HRDATA_S14
;
else
assign
CAHBLTIIO0I
=
32
'h
0
;
if
(
CAHBLTlIO0
[
15
]
)
assign
CAHBLTlIO0I
=
HRDATA_S15
;
else
assign
CAHBLTlIO0I
=
32
'h
0
;
if
(
CAHBLTlIO0
[
16
]
)
assign
CAHBLTOlO0I
=
HRDATA_S16
;
else
assign
CAHBLTOlO0I
=
32
'h
0
;
if
(
CAHBLTlIlll
[
0
]
)
assign
CAHBLTIIOl0
=
HRDATA_S0
;
else
assign
CAHBLTIIOl0
=
32
'h
0
;
if
(
CAHBLTlIlll
[
1
]
)
assign
CAHBLTlIOl0
=
HRDATA_S1
;
else
assign
CAHBLTlIOl0
=
32
'h
0
;
if
(
CAHBLTlIlll
[
2
]
)
assign
CAHBLTOlOl0
=
HRDATA_S2
;
else
assign
CAHBLTOlOl0
=
32
'h
0
;
if
(
CAHBLTlIlll
[
3
]
)
assign
CAHBLTIlOl0
=
HRDATA_S3
;
else
assign
CAHBLTIlOl0
=
32
'h
0
;
if
(
CAHBLTlIlll
[
4
]
)
assign
CAHBLTllOl0
=
HRDATA_S4
;
else
assign
CAHBLTllOl0
=
32
'h
0
;
if
(
CAHBLTlIlll
[
5
]
)
assign
CAHBLTO0Ol0
=
HRDATA_S5
;
else
assign
CAHBLTO0Ol0
=
32
'h
0
;
if
(
CAHBLTlIlll
[
6
]
)
assign
CAHBLTI0Ol0
=
HRDATA_S6
;
else
assign
CAHBLTI0Ol0
=
32
'h
0
;
if
(
CAHBLTlIlll
[
7
]
)
assign
CAHBLTl0Ol0
=
HRDATA_S7
;
else
assign
CAHBLTl0Ol0
=
32
'h
0
;
if
(
CAHBLTlIlll
[
8
]
)
assign
CAHBLTO1Ol0
=
HRDATA_S8
;
else
assign
CAHBLTO1Ol0
=
32
'h
0
;
if
(
CAHBLTlIlll
[
9
]
)
assign
CAHBLTI1Ol0
=
HRDATA_S9
;
else
assign
CAHBLTI1Ol0
=
32
'h
0
;
if
(
CAHBLTlIlll
[
10
]
)
assign
CAHBLTl1Ol0
=
HRDATA_S10
;
else
assign
CAHBLTl1Ol0
=
32
'h
0
;
if
(
CAHBLTlIlll
[
11
]
)
assign
CAHBLTOOIl0
=
HRDATA_S11
;
else
assign
CAHBLTOOIl0
=
32
'h
0
;
if
(
CAHBLTlIlll
[
12
]
)
assign
CAHBLTIOIl0
=
HRDATA_S12
;
else
assign
CAHBLTIOIl0
=
32
'h
0
;
if
(
CAHBLTlIlll
[
13
]
)
assign
CAHBLTlOIl0
=
HRDATA_S13
;
else
assign
CAHBLTlOIl0
=
32
'h
0
;
if
(
CAHBLTlIlll
[
14
]
)
assign
CAHBLTOIIl0
=
HRDATA_S14
;
else
assign
CAHBLTOIIl0
=
32
'h
0
;
if
(
CAHBLTlIlll
[
15
]
)
assign
CAHBLTIIIl0
=
HRDATA_S15
;
else
assign
CAHBLTIIIl0
=
32
'h
0
;
if
(
CAHBLTlIlll
[
16
]
)
assign
CAHBLTlIIl0
=
HRDATA_S16
;
else
assign
CAHBLTlIIl0
=
32
'h
0
;
if
(
CAHBLTOllll
[
0
]
)
assign
CAHBLTOlIl0
=
HRDATA_S0
;
else
assign
CAHBLTOlIl0
=
32
'h
0
;
if
(
CAHBLTOllll
[
1
]
)
assign
CAHBLTIlIl0
=
HRDATA_S1
;
else
assign
CAHBLTIlIl0
=
32
'h
0
;
if
(
CAHBLTOllll
[
2
]
)
assign
CAHBLTllIl0
=
HRDATA_S2
;
else
assign
CAHBLTllIl0
=
32
'h
0
;
if
(
CAHBLTOllll
[
3
]
)
assign
CAHBLTO0Il0
=
HRDATA_S3
;
else
assign
CAHBLTO0Il0
=
32
'h
0
;
if
(
CAHBLTOllll
[
4
]
)
assign
CAHBLTI0Il0
=
HRDATA_S4
;
else
assign
CAHBLTI0Il0
=
32
'h
0
;
if
(
CAHBLTOllll
[
5
]
)
assign
CAHBLTl0Il0
=
HRDATA_S5
;
else
assign
CAHBLTl0Il0
=
32
'h
0
;
if
(
CAHBLTOllll
[
6
]
)
assign
CAHBLTO1Il0
=
HRDATA_S6
;
else
assign
CAHBLTO1Il0
=
32
'h
0
;
if
(
CAHBLTOllll
[
7
]
)
assign
CAHBLTI1Il0
=
HRDATA_S7
;
else
assign
CAHBLTI1Il0
=
32
'h
0
;
if
(
CAHBLTOllll
[
8
]
)
assign
CAHBLTl1Il0
=
HRDATA_S8
;
else
assign
CAHBLTl1Il0
=
32
'h
0
;
if
(
CAHBLTOllll
[
9
]
)
assign
CAHBLTOOll0
=
HRDATA_S9
;
else
assign
CAHBLTOOll0
=
32
'h
0
;
if
(
CAHBLTOllll
[
10
]
)
assign
CAHBLTIOll0
=
HRDATA_S10
;
else
assign
CAHBLTIOll0
=
32
'h
0
;
if
(
CAHBLTOllll
[
11
]
)
assign
CAHBLTlOll0
=
HRDATA_S11
;
else
assign
CAHBLTlOll0
=
32
'h
0
;
if
(
CAHBLTOllll
[
12
]
)
assign
CAHBLTOIll0
=
HRDATA_S12
;
else
assign
CAHBLTOIll0
=
32
'h
0
;
if
(
CAHBLTOllll
[
13
]
)
assign
CAHBLTIIll0
=
HRDATA_S13
;
else
assign
CAHBLTIIll0
=
32
'h
0
;
if
(
CAHBLTOllll
[
14
]
)
assign
CAHBLTlIll0
=
HRDATA_S14
;
else
assign
CAHBLTlIll0
=
32
'h
0
;
if
(
CAHBLTOllll
[
15
]
)
assign
CAHBLTOlll0
=
HRDATA_S15
;
else
assign
CAHBLTOlll0
=
32
'h
0
;
if
(
CAHBLTOllll
[
16
]
)
assign
CAHBLTIlll0
=
HRDATA_S16
;
else
assign
CAHBLTIlll0
=
32
'h
0
;
endgenerate
generate
if
(
CAHBLTIIO0
[
0
]
)
assign
CAHBLTOOO1I
=
HWDATA_M0
;
else
assign
CAHBLTOOO1I
=
32
'h
0
;
if
(
CAHBLTIIO0
[
1
]
)
assign
CAHBLTIOO1I
=
HWDATA_M0
;
else
assign
CAHBLTIOO1I
=
32
'h
0
;
if
(
CAHBLTIIO0
[
2
]
)
assign
CAHBLTlOO1I
=
HWDATA_M0
;
else
assign
CAHBLTlOO1I
=
32
'h
0
;
if
(
CAHBLTIIO0
[
3
]
)
assign
CAHBLTOIO1I
=
HWDATA_M0
;
else
assign
CAHBLTOIO1I
=
32
'h
0
;
if
(
CAHBLTIIO0
[
4
]
)
assign
CAHBLTIIO1I
=
HWDATA_M0
;
else
assign
CAHBLTIIO1I
=
32
'h
0
;
if
(
CAHBLTIIO0
[
5
]
)
assign
CAHBLTlIO1I
=
HWDATA_M0
;
else
assign
CAHBLTlIO1I
=
32
'h
0
;
if
(
CAHBLTIIO0
[
6
]
)
assign
CAHBLTOlO1I
=
HWDATA_M0
;
else
assign
CAHBLTOlO1I
=
32
'h
0
;
if
(
CAHBLTIIO0
[
7
]
)
assign
CAHBLTIlO1I
=
HWDATA_M0
;
else
assign
CAHBLTIlO1I
=
32
'h
0
;
if
(
CAHBLTIIO0
[
8
]
)
assign
CAHBLTllO1I
=
HWDATA_M0
;
else
assign
CAHBLTllO1I
=
32
'h
0
;
if
(
CAHBLTIIO0
[
9
]
)
assign
CAHBLTO0O1I
=
HWDATA_M0
;
else
assign
CAHBLTO0O1I
=
32
'h
0
;
if
(
CAHBLTIIO0
[
10
]
)
assign
CAHBLTI0O1I
=
HWDATA_M0
;
else
assign
CAHBLTI0O1I
=
32
'h
0
;
if
(
CAHBLTIIO0
[
11
]
)
assign
CAHBLTl0O1I
=
HWDATA_M0
;
else
assign
CAHBLTl0O1I
=
32
'h
0
;
if
(
CAHBLTIIO0
[
12
]
)
assign
CAHBLTO1O1I
=
HWDATA_M0
;
else
assign
CAHBLTO1O1I
=
32
'h
0
;
if
(
CAHBLTIIO0
[
13
]
)
assign
CAHBLTI1O1I
=
HWDATA_M0
;
else
assign
CAHBLTI1O1I
=
32
'h
0
;
if
(
CAHBLTIIO0
[
14
]
)
assign
CAHBLTl1O1I
=
HWDATA_M0
;
else
assign
CAHBLTl1O1I
=
32
'h
0
;
if
(
CAHBLTIIO0
[
15
]
)
assign
CAHBLTOOI1I
=
HWDATA_M0
;
else
assign
CAHBLTOOI1I
=
32
'h
0
;
if
(
CAHBLTIIO0
[
16
]
)
assign
CAHBLTIOI1I
=
HWDATA_M0
;
else
assign
CAHBLTIOI1I
=
32
'h
0
;
if
(
CAHBLTlIO0
[
0
]
)
assign
CAHBLTlOI1I
=
HWDATA_M1
;
else
assign
CAHBLTlOI1I
=
32
'h
0
;
if
(
CAHBLTlIO0
[
1
]
)
assign
CAHBLTOII1I
=
HWDATA_M1
;
else
assign
CAHBLTOII1I
=
32
'h
0
;
if
(
CAHBLTlIO0
[
2
]
)
assign
CAHBLTIII1I
=
HWDATA_M1
;
else
assign
CAHBLTIII1I
=
32
'h
0
;
if
(
CAHBLTlIO0
[
3
]
)
assign
CAHBLTlII1I
=
HWDATA_M1
;
else
assign
CAHBLTlII1I
=
32
'h
0
;
if
(
CAHBLTlIO0
[
4
]
)
assign
CAHBLTOlI1I
=
HWDATA_M1
;
else
assign
CAHBLTOlI1I
=
32
'h
0
;
if
(
CAHBLTlIO0
[
5
]
)
assign
CAHBLTIlI1I
=
HWDATA_M1
;
else
assign
CAHBLTIlI1I
=
32
'h
0
;
if
(
CAHBLTlIO0
[
6
]
)
assign
CAHBLTllI1I
=
HWDATA_M1
;
else
assign
CAHBLTllI1I
=
32
'h
0
;
if
(
CAHBLTlIO0
[
7
]
)
assign
CAHBLTO0I1I
=
HWDATA_M1
;
else
assign
CAHBLTO0I1I
=
32
'h
0
;
if
(
CAHBLTlIO0
[
8
]
)
assign
CAHBLTI0I1I
=
HWDATA_M1
;
else
assign
CAHBLTI0I1I
=
32
'h
0
;
if
(
CAHBLTlIO0
[
9
]
)
assign
CAHBLTl0I1I
=
HWDATA_M1
;
else
assign
CAHBLTl0I1I
=
32
'h
0
;
if
(
CAHBLTlIO0
[
10
]
)
assign
CAHBLTO1I1I
=
HWDATA_M1
;
else
assign
CAHBLTO1I1I
=
32
'h
0
;
if
(
CAHBLTlIO0
[
11
]
)
assign
CAHBLTI1I1I
=
HWDATA_M1
;
else
assign
CAHBLTI1I1I
=
32
'h
0
;
if
(
CAHBLTlIO0
[
12
]
)
assign
CAHBLTl1I1I
=
HWDATA_M1
;
else
assign
CAHBLTl1I1I
=
32
'h
0
;
if
(
CAHBLTlIO0
[
13
]
)
assign
CAHBLTOOl1I
=
HWDATA_M1
;
else
assign
CAHBLTOOl1I
=
32
'h
0
;
if
(
CAHBLTlIO0
[
14
]
)
assign
CAHBLTIOl1I
=
HWDATA_M1
;
else
assign
CAHBLTIOl1I
=
32
'h
0
;
if
(
CAHBLTlIO0
[
15
]
)
assign
CAHBLTlOl1I
=
HWDATA_M1
;
else
assign
CAHBLTlOl1I
=
32
'h
0
;
if
(
CAHBLTlIO0
[
16
]
)
assign
CAHBLTOIl1I
=
HWDATA_M1
;
else
assign
CAHBLTOIl1I
=
32
'h
0
;
if
(
CAHBLTlIlll
[
0
]
)
assign
CAHBLTO11l0
=
HWDATA_M2
;
else
assign
CAHBLTO11l0
=
32
'h
0
;
if
(
CAHBLTlIlll
[
1
]
)
assign
CAHBLTI11l0
=
HWDATA_M2
;
else
assign
CAHBLTI11l0
=
32
'h
0
;
if
(
CAHBLTlIlll
[
2
]
)
assign
CAHBLTl11l0
=
HWDATA_M2
;
else
assign
CAHBLTl11l0
=
32
'h
0
;
if
(
CAHBLTlIlll
[
3
]
)
assign
CAHBLTOOO00
=
HWDATA_M2
;
else
assign
CAHBLTOOO00
=
32
'h
0
;
if
(
CAHBLTlIlll
[
4
]
)
assign
CAHBLTIOO00
=
HWDATA_M2
;
else
assign
CAHBLTIOO00
=
32
'h
0
;
if
(
CAHBLTlIlll
[
5
]
)
assign
CAHBLTlOO00
=
HWDATA_M2
;
else
assign
CAHBLTlOO00
=
32
'h
0
;
if
(
CAHBLTlIlll
[
6
]
)
assign
CAHBLTOIO00
=
HWDATA_M2
;
else
assign
CAHBLTOIO00
=
32
'h
0
;
if
(
CAHBLTlIlll
[
7
]
)
assign
CAHBLTIIO00
=
HWDATA_M2
;
else
assign
CAHBLTIIO00
=
32
'h
0
;
if
(
CAHBLTlIlll
[
8
]
)
assign
CAHBLTlIO00
=
HWDATA_M2
;
else
assign
CAHBLTlIO00
=
32
'h
0
;
if
(
CAHBLTlIlll
[
9
]
)
assign
CAHBLTOlO00
=
HWDATA_M2
;
else
assign
CAHBLTOlO00
=
32
'h
0
;
if
(
CAHBLTlIlll
[
10
]
)
assign
CAHBLTIlO00
=
HWDATA_M2
;
else
assign
CAHBLTIlO00
=
32
'h
0
;
if
(
CAHBLTlIlll
[
11
]
)
assign
CAHBLTllO00
=
HWDATA_M2
;
else
assign
CAHBLTllO00
=
32
'h
0
;
if
(
CAHBLTlIlll
[
12
]
)
assign
CAHBLTO0O00
=
HWDATA_M2
;
else
assign
CAHBLTO0O00
=
32
'h
0
;
if
(
CAHBLTlIlll
[
13
]
)
assign
CAHBLTI0O00
=
HWDATA_M2
;
else
assign
CAHBLTI0O00
=
32
'h
0
;
if
(
CAHBLTlIlll
[
14
]
)
assign
CAHBLTl0O00
=
HWDATA_M2
;
else
assign
CAHBLTl0O00
=
32
'h
0
;
if
(
CAHBLTlIlll
[
15
]
)
assign
CAHBLTO1O00
=
HWDATA_M2
;
else
assign
CAHBLTO1O00
=
32
'h
0
;
if
(
CAHBLTlIlll
[
16
]
)
assign
CAHBLTI1O00
=
HWDATA_M2
;
else
assign
CAHBLTI1O00
=
32
'h
0
;
if
(
CAHBLTOllll
[
0
]
)
assign
CAHBLTl1O00
=
HWDATA_M3
;
else
assign
CAHBLTl1O00
=
32
'h
0
;
if
(
CAHBLTOllll
[
1
]
)
assign
CAHBLTOOI00
=
HWDATA_M3
;
else
assign
CAHBLTOOI00
=
32
'h
0
;
if
(
CAHBLTOllll
[
2
]
)
assign
CAHBLTIOI00
=
HWDATA_M3
;
else
assign
CAHBLTIOI00
=
32
'h
0
;
if
(
CAHBLTOllll
[
3
]
)
assign
CAHBLTlOI00
=
HWDATA_M3
;
else
assign
CAHBLTlOI00
=
32
'h
0
;
if
(
CAHBLTOllll
[
4
]
)
assign
CAHBLTOII00
=
HWDATA_M3
;
else
assign
CAHBLTOII00
=
32
'h
0
;
if
(
CAHBLTOllll
[
5
]
)
assign
CAHBLTIII00
=
HWDATA_M3
;
else
assign
CAHBLTIII00
=
32
'h
0
;
if
(
CAHBLTOllll
[
6
]
)
assign
CAHBLTlII00
=
HWDATA_M3
;
else
assign
CAHBLTlII00
=
32
'h
0
;
if
(
CAHBLTOllll
[
7
]
)
assign
CAHBLTOlI00
=
HWDATA_M3
;
else
assign
CAHBLTOlI00
=
32
'h
0
;
if
(
CAHBLTOllll
[
8
]
)
assign
CAHBLTIlI00
=
HWDATA_M3
;
else
assign
CAHBLTIlI00
=
32
'h
0
;
if
(
CAHBLTOllll
[
9
]
)
assign
CAHBLTllI00
=
HWDATA_M3
;
else
assign
CAHBLTllI00
=
32
'h
0
;
if
(
CAHBLTOllll
[
10
]
)
assign
CAHBLTO0I00
=
HWDATA_M3
;
else
assign
CAHBLTO0I00
=
32
'h
0
;
if
(
CAHBLTOllll
[
11
]
)
assign
CAHBLTI0I00
=
HWDATA_M3
;
else
assign
CAHBLTI0I00
=
32
'h
0
;
if
(
CAHBLTOllll
[
12
]
)
assign
CAHBLTl0I00
=
HWDATA_M3
;
else
assign
CAHBLTl0I00
=
32
'h
0
;
if
(
CAHBLTOllll
[
13
]
)
assign
CAHBLTO1I00
=
HWDATA_M3
;
else
assign
CAHBLTO1I00
=
32
'h
0
;
if
(
CAHBLTOllll
[
14
]
)
assign
CAHBLTI1I00
=
HWDATA_M3
;
else
assign
CAHBLTI1I00
=
32
'h
0
;
if
(
CAHBLTOllll
[
15
]
)
assign
CAHBLTl1I00
=
HWDATA_M3
;
else
assign
CAHBLTl1I00
=
32
'h
0
;
if
(
CAHBLTOllll
[
16
]
)
assign
CAHBLTOOl00
=
HWDATA_M3
;
else
assign
CAHBLTOOl00
=
32
'h
0
;
endgenerate
generate
if
(
CAHBLTIIO0
[
0
]
)
assign
CAHBLTIlO0I
=
HREADYOUT_S0
;
else
assign
CAHBLTIlO0I
=
1
'b
1
;
if
(
CAHBLTIIO0
[
1
]
)
assign
CAHBLTllO0I
=
HREADYOUT_S1
;
else
assign
CAHBLTllO0I
=
1
'b
1
;
if
(
CAHBLTIIO0
[
2
]
)
assign
CAHBLTO0O0I
=
HREADYOUT_S2
;
else
assign
CAHBLTO0O0I
=
1
'b
1
;
if
(
CAHBLTIIO0
[
3
]
)
assign
CAHBLTI0O0I
=
HREADYOUT_S3
;
else
assign
CAHBLTI0O0I
=
1
'b
1
;
if
(
CAHBLTIIO0
[
4
]
)
assign
CAHBLTl0O0I
=
HREADYOUT_S4
;
else
assign
CAHBLTl0O0I
=
1
'b
1
;
if
(
CAHBLTIIO0
[
5
]
)
assign
CAHBLTO1O0I
=
HREADYOUT_S5
;
else
assign
CAHBLTO1O0I
=
1
'b
1
;
if
(
CAHBLTIIO0
[
6
]
)
assign
CAHBLTI1O0I
=
HREADYOUT_S6
;
else
assign
CAHBLTI1O0I
=
1
'b
1
;
if
(
CAHBLTIIO0
[
7
]
)
assign
CAHBLTl1O0I
=
HREADYOUT_S7
;
else
assign
CAHBLTl1O0I
=
1
'b
1
;
if
(
CAHBLTIIO0
[
8
]
)
assign
CAHBLTOOI0I
=
HREADYOUT_S8
;
else
assign
CAHBLTOOI0I
=
1
'b
1
;
if
(
CAHBLTIIO0
[
9
]
)
assign
CAHBLTIOI0I
=
HREADYOUT_S9
;
else
assign
CAHBLTIOI0I
=
1
'b
1
;
if
(
CAHBLTIIO0
[
10
]
)
assign
CAHBLTlOI0I
=
HREADYOUT_S10
;
else
assign
CAHBLTlOI0I
=
1
'b
1
;
if
(
CAHBLTIIO0
[
11
]
)
assign
CAHBLTOII0I
=
HREADYOUT_S11
;
else
assign
CAHBLTOII0I
=
1
'b
1
;
if
(
CAHBLTIIO0
[
12
]
)
assign
CAHBLTIII0I
=
HREADYOUT_S12
;
else
assign
CAHBLTIII0I
=
1
'b
1
;
if
(
CAHBLTIIO0
[
13
]
)
assign
CAHBLTlII0I
=
HREADYOUT_S13
;
else
assign
CAHBLTlII0I
=
1
'b
1
;
if
(
CAHBLTIIO0
[
14
]
)
assign
CAHBLTOlI0I
=
HREADYOUT_S14
;
else
assign
CAHBLTOlI0I
=
1
'b
1
;
if
(
CAHBLTIIO0
[
15
]
)
assign
CAHBLTIlI0I
=
HREADYOUT_S15
;
else
assign
CAHBLTIlI0I
=
1
'b
1
;
if
(
CAHBLTIIO0
[
16
]
)
assign
CAHBLTllI0I
=
HREADYOUT_S16
;
else
assign
CAHBLTllI0I
=
1
'b
1
;
if
(
CAHBLTlIO0
[
0
]
)
assign
CAHBLTO0I0I
=
HREADYOUT_S0
;
else
assign
CAHBLTO0I0I
=
1
'b
1
;
if
(
CAHBLTlIO0
[
1
]
)
assign
CAHBLTI0I0I
=
HREADYOUT_S1
;
else
assign
CAHBLTI0I0I
=
1
'b
1
;
if
(
CAHBLTlIO0
[
2
]
)
assign
CAHBLTl0I0I
=
HREADYOUT_S2
;
else
assign
CAHBLTl0I0I
=
1
'b
1
;
if
(
CAHBLTlIO0
[
3
]
)
assign
CAHBLTO1I0I
=
HREADYOUT_S3
;
else
assign
CAHBLTO1I0I
=
1
'b
1
;
if
(
CAHBLTlIO0
[
4
]
)
assign
CAHBLTI1I0I
=
HREADYOUT_S4
;
else
assign
CAHBLTI1I0I
=
1
'b
1
;
if
(
CAHBLTlIO0
[
5
]
)
assign
CAHBLTl1I0I
=
HREADYOUT_S5
;
else
assign
CAHBLTl1I0I
=
1
'b
1
;
if
(
CAHBLTlIO0
[
6
]
)
assign
CAHBLTOOl0I
=
HREADYOUT_S6
;
else
assign
CAHBLTOOl0I
=
1
'b
1
;
if
(
CAHBLTlIO0
[
7
]
)
assign
CAHBLTIOl0I
=
HREADYOUT_S7
;
else
assign
CAHBLTIOl0I
=
1
'b
1
;
if
(
CAHBLTlIO0
[
8
]
)
assign
CAHBLTlOl0I
=
HREADYOUT_S8
;
else
assign
CAHBLTlOl0I
=
1
'b
1
;
if
(
CAHBLTlIO0
[
9
]
)
assign
CAHBLTOIl0I
=
HREADYOUT_S9
;
else
assign
CAHBLTOIl0I
=
1
'b
1
;
if
(
CAHBLTlIO0
[
10
]
)
assign
CAHBLTIIl0I
=
HREADYOUT_S10
;
else
assign
CAHBLTIIl0I
=
1
'b
1
;
if
(
CAHBLTlIO0
[
11
]
)
assign
CAHBLTlIl0I
=
HREADYOUT_S11
;
else
assign
CAHBLTlIl0I
=
1
'b
1
;
if
(
CAHBLTlIO0
[
12
]
)
assign
CAHBLTOll0I
=
HREADYOUT_S12
;
else
assign
CAHBLTOll0I
=
1
'b
1
;
if
(
CAHBLTlIO0
[
13
]
)
assign
CAHBLTIll0I
=
HREADYOUT_S13
;
else
assign
CAHBLTIll0I
=
1
'b
1
;
if
(
CAHBLTlIO0
[
14
]
)
assign
CAHBLTlll0I
=
HREADYOUT_S14
;
else
assign
CAHBLTlll0I
=
1
'b
1
;
if
(
CAHBLTlIO0
[
15
]
)
assign
CAHBLTO0l0I
=
HREADYOUT_S15
;
else
assign
CAHBLTO0l0I
=
1
'b
1
;
if
(
CAHBLTlIO0
[
16
]
)
assign
CAHBLTI0l0I
=
HREADYOUT_S16
;
else
assign
CAHBLTI0l0I
=
1
'b
1
;
if
(
CAHBLTlIlll
[
0
]
)
assign
CAHBLTllll0
=
HREADYOUT_S0
;
else
assign
CAHBLTllll0
=
1
'b
1
;
if
(
CAHBLTlIlll
[
1
]
)
assign
CAHBLTO0ll0
=
HREADYOUT_S1
;
else
assign
CAHBLTO0ll0
=
1
'b
1
;
if
(
CAHBLTlIlll
[
2
]
)
assign
CAHBLTI0ll0
=
HREADYOUT_S2
;
else
assign
CAHBLTI0ll0
=
1
'b
1
;
if
(
CAHBLTlIlll
[
3
]
)
assign
CAHBLTl0ll0
=
HREADYOUT_S3
;
else
assign
CAHBLTl0ll0
=
1
'b
1
;
if
(
CAHBLTlIlll
[
4
]
)
assign
CAHBLTO1ll0
=
HREADYOUT_S4
;
else
assign
CAHBLTO1ll0
=
1
'b
1
;
if
(
CAHBLTlIlll
[
5
]
)
assign
CAHBLTI1ll0
=
HREADYOUT_S5
;
else
assign
CAHBLTI1ll0
=
1
'b
1
;
if
(
CAHBLTlIlll
[
6
]
)
assign
CAHBLTl1ll0
=
HREADYOUT_S6
;
else
assign
CAHBLTl1ll0
=
1
'b
1
;
if
(
CAHBLTlIlll
[
7
]
)
assign
CAHBLTOO0l0
=
HREADYOUT_S7
;
else
assign
CAHBLTOO0l0
=
1
'b
1
;
if
(
CAHBLTlIlll
[
8
]
)
assign
CAHBLTIO0l0
=
HREADYOUT_S8
;
else
assign
CAHBLTIO0l0
=
1
'b
1
;
if
(
CAHBLTlIlll
[
9
]
)
assign
CAHBLTlO0l0
=
HREADYOUT_S9
;
else
assign
CAHBLTlO0l0
=
1
'b
1
;
if
(
CAHBLTlIlll
[
10
]
)
assign
CAHBLTOI0l0
=
HREADYOUT_S10
;
else
assign
CAHBLTOI0l0
=
1
'b
1
;
if
(
CAHBLTlIlll
[
11
]
)
assign
CAHBLTII0l0
=
HREADYOUT_S11
;
else
assign
CAHBLTII0l0
=
1
'b
1
;
if
(
CAHBLTlIlll
[
12
]
)
assign
CAHBLTlI0l0
=
HREADYOUT_S12
;
else
assign
CAHBLTlI0l0
=
1
'b
1
;
if
(
CAHBLTlIlll
[
13
]
)
assign
CAHBLTOl0l0
=
HREADYOUT_S13
;
else
assign
CAHBLTOl0l0
=
1
'b
1
;
if
(
CAHBLTlIlll
[
14
]
)
assign
CAHBLTIl0l0
=
HREADYOUT_S14
;
else
assign
CAHBLTIl0l0
=
1
'b
1
;
if
(
CAHBLTlIlll
[
15
]
)
assign
CAHBLTll0l0
=
HREADYOUT_S15
;
else
assign
CAHBLTll0l0
=
1
'b
1
;
if
(
CAHBLTlIlll
[
16
]
)
assign
CAHBLTO00l0
=
HREADYOUT_S16
;
else
assign
CAHBLTO00l0
=
1
'b
1
;
if
(
CAHBLTOllll
[
0
]
)
assign
CAHBLTI00l0
=
HREADYOUT_S0
;
else
assign
CAHBLTI00l0
=
1
'b
1
;
if
(
CAHBLTOllll
[
1
]
)
assign
CAHBLTl00l0
=
HREADYOUT_S1
;
else
assign
CAHBLTl00l0
=
1
'b
1
;
if
(
CAHBLTOllll
[
2
]
)
assign
CAHBLTO10l0
=
HREADYOUT_S2
;
else
assign
CAHBLTO10l0
=
1
'b
1
;
if
(
CAHBLTOllll
[
3
]
)
assign
CAHBLTI10l0
=
HREADYOUT_S3
;
else
assign
CAHBLTI10l0
=
1
'b
1
;
if
(
CAHBLTOllll
[
4
]
)
assign
CAHBLTl10l0
=
HREADYOUT_S4
;
else
assign
CAHBLTl10l0
=
1
'b
1
;
if
(
CAHBLTOllll
[
5
]
)
assign
CAHBLTOO1l0
=
HREADYOUT_S5
;
else
assign
CAHBLTOO1l0
=
1
'b
1
;
if
(
CAHBLTOllll
[
6
]
)
assign
CAHBLTIO1l0
=
HREADYOUT_S6
;
else
assign
CAHBLTIO1l0
=
1
'b
1
;
if
(
CAHBLTOllll
[
7
]
)
assign
CAHBLTlO1l0
=
HREADYOUT_S7
;
else
assign
CAHBLTlO1l0
=
1
'b
1
;
if
(
CAHBLTOllll
[
8
]
)
assign
CAHBLTOI1l0
=
HREADYOUT_S8
;
else
assign
CAHBLTOI1l0
=
1
'b
1
;
if
(
CAHBLTOllll
[
9
]
)
assign
CAHBLTII1l0
=
HREADYOUT_S9
;
else
assign
CAHBLTII1l0
=
1
'b
1
;
if
(
CAHBLTOllll
[
10
]
)
assign
CAHBLTlI1l0
=
HREADYOUT_S10
;
else
assign
CAHBLTlI1l0
=
1
'b
1
;
if
(
CAHBLTOllll
[
11
]
)
assign
CAHBLTOl1l0
=
HREADYOUT_S11
;
else
assign
CAHBLTOl1l0
=
1
'b
1
;
if
(
CAHBLTOllll
[
12
]
)
assign
CAHBLTIl1l0
=
HREADYOUT_S12
;
else
assign
CAHBLTIl1l0
=
1
'b
1
;
if
(
CAHBLTOllll
[
13
]
)
assign
CAHBLTll1l0
=
HREADYOUT_S13
;
else
assign
CAHBLTll1l0
=
1
'b
1
;
if
(
CAHBLTOllll
[
14
]
)
assign
CAHBLTO01l0
=
HREADYOUT_S14
;
else
assign
CAHBLTO01l0
=
1
'b
1
;
if
(
CAHBLTOllll
[
15
]
)
assign
CAHBLTI01l0
=
HREADYOUT_S15
;
else
assign
CAHBLTI01l0
=
1
'b
1
;
if
(
CAHBLTOllll
[
16
]
)
assign
CAHBLTl01l0
=
HREADYOUT_S16
;
else
assign
CAHBLTl01l0
=
1
'b
1
;
endgenerate
generate
if
(
CAHBLTIIO0
[
0
]
|
CAHBLTlIO0
[
0
]
|
CAHBLTlIlll
[
0
]
|
CAHBLTOllll
[
0
]
)
assign
CAHBLTl0l0I
=
HREADYOUT_S0
;
else
assign
CAHBLTl0l0I
=
1
'b
1
;
if
(
CAHBLTIIO0
[
1
]
|
CAHBLTlIO0
[
1
]
|
CAHBLTlIlll
[
1
]
|
CAHBLTOllll
[
1
]
)
assign
CAHBLTO1l0I
=
HREADYOUT_S1
;
else
assign
CAHBLTO1l0I
=
1
'b
1
;
if
(
CAHBLTIIO0
[
2
]
|
CAHBLTlIO0
[
2
]
|
CAHBLTlIlll
[
2
]
|
CAHBLTOllll
[
2
]
)
assign
CAHBLTI1l0I
=
HREADYOUT_S2
;
else
assign
CAHBLTI1l0I
=
1
'b
1
;
if
(
CAHBLTIIO0
[
3
]
|
CAHBLTlIO0
[
3
]
|
CAHBLTlIlll
[
3
]
|
CAHBLTOllll
[
3
]
)
assign
CAHBLTl1l0I
=
HREADYOUT_S3
;
else
assign
CAHBLTl1l0I
=
1
'b
1
;
if
(
CAHBLTIIO0
[
4
]
|
CAHBLTlIO0
[
4
]
|
CAHBLTlIlll
[
4
]
|
CAHBLTOllll
[
4
]
)
assign
CAHBLTOO00I
=
HREADYOUT_S4
;
else
assign
CAHBLTOO00I
=
1
'b
1
;
if
(
CAHBLTIIO0
[
5
]
|
CAHBLTlIO0
[
5
]
|
CAHBLTlIlll
[
5
]
|
CAHBLTOllll
[
5
]
)
assign
CAHBLTIO00I
=
HREADYOUT_S5
;
else
assign
CAHBLTIO00I
=
1
'b
1
;
if
(
CAHBLTIIO0
[
6
]
|
CAHBLTlIO0
[
6
]
|
CAHBLTlIlll
[
6
]
|
CAHBLTOllll
[
6
]
)
assign
CAHBLTlO00I
=
HREADYOUT_S6
;
else
assign
CAHBLTlO00I
=
1
'b
1
;
if
(
CAHBLTIIO0
[
7
]
|
CAHBLTlIO0
[
7
]
|
CAHBLTlIlll
[
7
]
|
CAHBLTOllll
[
7
]
)
assign
CAHBLTOI00I
=
HREADYOUT_S7
;
else
assign
CAHBLTOI00I
=
1
'b
1
;
if
(
CAHBLTIIO0
[
8
]
|
CAHBLTlIO0
[
8
]
|
CAHBLTlIlll
[
8
]
|
CAHBLTOllll
[
8
]
)
assign
CAHBLTII00I
=
HREADYOUT_S8
;
else
assign
CAHBLTII00I
=
1
'b
1
;
if
(
CAHBLTIIO0
[
9
]
|
CAHBLTlIO0
[
9
]
|
CAHBLTlIlll
[
9
]
|
CAHBLTOllll
[
9
]
)
assign
CAHBLTlI00I
=
HREADYOUT_S9
;
else
assign
CAHBLTlI00I
=
1
'b
1
;
if
(
CAHBLTIIO0
[
10
]
|
CAHBLTlIO0
[
10
]
|
CAHBLTlIlll
[
10
]
|
CAHBLTOllll
[
10
]
)
assign
CAHBLTOl00I
=
HREADYOUT_S10
;
else
assign
CAHBLTOl00I
=
1
'b
1
;
if
(
CAHBLTIIO0
[
11
]
|
CAHBLTlIO0
[
11
]
|
CAHBLTlIlll
[
11
]
|
CAHBLTOllll
[
11
]
)
assign
CAHBLTIl00I
=
HREADYOUT_S11
;
else
assign
CAHBLTIl00I
=
1
'b
1
;
if
(
CAHBLTIIO0
[
12
]
|
CAHBLTlIO0
[
12
]
|
CAHBLTlIlll
[
12
]
|
CAHBLTOllll
[
12
]
)
assign
CAHBLTll00I
=
HREADYOUT_S12
;
else
assign
CAHBLTll00I
=
1
'b
1
;
if
(
CAHBLTIIO0
[
13
]
|
CAHBLTlIO0
[
13
]
|
CAHBLTlIlll
[
13
]
|
CAHBLTOllll
[
13
]
)
assign
CAHBLTO000I
=
HREADYOUT_S13
;
else
assign
CAHBLTO000I
=
1
'b
1
;
if
(
CAHBLTIIO0
[
14
]
|
CAHBLTlIO0
[
14
]
|
CAHBLTlIlll
[
14
]
|
CAHBLTOllll
[
14
]
)
assign
CAHBLTI000I
=
HREADYOUT_S14
;
else
assign
CAHBLTI000I
=
1
'b
1
;
if
(
CAHBLTIIO0
[
15
]
|
CAHBLTlIO0
[
15
]
|
CAHBLTlIlll
[
15
]
|
CAHBLTOllll
[
15
]
)
assign
CAHBLTl000I
=
HREADYOUT_S15
;
else
assign
CAHBLTl000I
=
1
'b
1
;
if
(
CAHBLTIIO0
[
16
]
|
CAHBLTlIO0
[
16
]
|
CAHBLTlIlll
[
16
]
|
CAHBLTOllll
[
16
]
)
assign
CAHBLTO100I
=
HREADYOUT_S16
;
else
assign
CAHBLTO100I
=
1
'b
1
;
endgenerate
generate
if
(
CAHBLTIIO0
[
0
]
|
CAHBLTlIO0
[
0
]
|
CAHBLTlIlll
[
0
]
|
CAHBLTOllll
[
0
]
)
assign
CAHBLTI100I
=
HRESP_S0
;
else
assign
CAHBLTI100I
=
1
'b
0
;
if
(
CAHBLTIIO0
[
1
]
|
CAHBLTlIO0
[
1
]
|
CAHBLTlIlll
[
1
]
|
CAHBLTOllll
[
1
]
)
assign
CAHBLTl100I
=
HRESP_S1
;
else
assign
CAHBLTl100I
=
1
'b
0
;
if
(
CAHBLTIIO0
[
2
]
|
CAHBLTlIO0
[
2
]
|
CAHBLTlIlll
[
2
]
|
CAHBLTOllll
[
2
]
)
assign
CAHBLTOO10I
=
HRESP_S2
;
else
assign
CAHBLTOO10I
=
1
'b
0
;
if
(
CAHBLTIIO0
[
3
]
|
CAHBLTlIO0
[
3
]
|
CAHBLTlIlll
[
3
]
|
CAHBLTOllll
[
3
]
)
assign
CAHBLTIO10I
=
HRESP_S3
;
else
assign
CAHBLTIO10I
=
1
'b
0
;
if
(
CAHBLTIIO0
[
4
]
|
CAHBLTlIO0
[
4
]
|
CAHBLTlIlll
[
4
]
|
CAHBLTOllll
[
4
]
)
assign
CAHBLTlO10I
=
HRESP_S4
;
else
assign
CAHBLTlO10I
=
1
'b
0
;
if
(
CAHBLTIIO0
[
5
]
|
CAHBLTlIO0
[
5
]
|
CAHBLTlIlll
[
5
]
|
CAHBLTOllll
[
5
]
)
assign
CAHBLTOI10I
=
HRESP_S5
;
else
assign
CAHBLTOI10I
=
1
'b
0
;
if
(
CAHBLTIIO0
[
6
]
|
CAHBLTlIO0
[
6
]
|
CAHBLTlIlll
[
6
]
|
CAHBLTOllll
[
6
]
)
assign
CAHBLTII10I
=
HRESP_S6
;
else
assign
CAHBLTII10I
=
1
'b
0
;
if
(
CAHBLTIIO0
[
7
]
|
CAHBLTlIO0
[
7
]
|
CAHBLTlIlll
[
7
]
|
CAHBLTOllll
[
7
]
)
assign
CAHBLTlI10I
=
HRESP_S7
;
else
assign
CAHBLTlI10I
=
1
'b
0
;
if
(
CAHBLTIIO0
[
8
]
|
CAHBLTlIO0
[
8
]
|
CAHBLTlIlll
[
8
]
|
CAHBLTOllll
[
8
]
)
assign
CAHBLTOl10I
=
HRESP_S8
;
else
assign
CAHBLTOl10I
=
1
'b
0
;
if
(
CAHBLTIIO0
[
9
]
|
CAHBLTlIO0
[
9
]
|
CAHBLTlIlll
[
9
]
|
CAHBLTOllll
[
9
]
)
assign
CAHBLTIl10I
=
HRESP_S9
;
else
assign
CAHBLTIl10I
=
1
'b
0
;
if
(
CAHBLTIIO0
[
10
]
|
CAHBLTlIO0
[
10
]
|
CAHBLTlIlll
[
10
]
|
CAHBLTOllll
[
10
]
)
assign
CAHBLTll10I
=
HRESP_S10
;
else
assign
CAHBLTll10I
=
1
'b
0
;
if
(
CAHBLTIIO0
[
11
]
|
CAHBLTlIO0
[
11
]
|
CAHBLTlIlll
[
11
]
|
CAHBLTOllll
[
11
]
)
assign
CAHBLTO010I
=
HRESP_S11
;
else
assign
CAHBLTO010I
=
1
'b
0
;
if
(
CAHBLTIIO0
[
12
]
|
CAHBLTlIO0
[
12
]
|
CAHBLTlIlll
[
12
]
|
CAHBLTOllll
[
12
]
)
assign
CAHBLTI010I
=
HRESP_S12
;
else
assign
CAHBLTI010I
=
1
'b
0
;
if
(
CAHBLTIIO0
[
13
]
|
CAHBLTlIO0
[
13
]
|
CAHBLTlIlll
[
13
]
|
CAHBLTOllll
[
13
]
)
assign
CAHBLTl010I
=
HRESP_S13
;
else
assign
CAHBLTl010I
=
1
'b
0
;
if
(
CAHBLTIIO0
[
14
]
|
CAHBLTlIO0
[
14
]
|
CAHBLTlIlll
[
14
]
|
CAHBLTOllll
[
14
]
)
assign
CAHBLTO110I
=
HRESP_S14
;
else
assign
CAHBLTO110I
=
1
'b
0
;
if
(
CAHBLTIIO0
[
15
]
|
CAHBLTlIO0
[
15
]
|
CAHBLTlIlll
[
15
]
|
CAHBLTOllll
[
15
]
)
assign
CAHBLTI110I
=
HRESP_S15
;
else
assign
CAHBLTI110I
=
1
'b
0
;
if
(
CAHBLTIIO0
[
16
]
|
CAHBLTlIO0
[
16
]
|
CAHBLTlIlll
[
16
]
|
CAHBLTOllll
[
16
]
)
assign
CAHBLTl110I
=
HRESP_S16
;
else
assign
CAHBLTl110I
=
1
'b
0
;
endgenerate
CAHBLTIIOI
#
(
.MEMSPACE
(
MEMSPACE
)
,
.HADDR_SHG_CFG
(
HADDR_SHG_CFG
)
,
.CAHBLTI
(
CAHBLTI
)
,
.CAHBLTl
(
CAHBLTIIO0
)
,
.SYNC_RESET
(
SYNC_RESET
)
)
CAHBLTOOIll
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.CAHBLTlIOI
(
HADDR_M0
)
,
.CAHBLTOlOI
(
HMASTLOCK_M0
)
,
.CAHBLTIlOI
(
HSIZE_M0
)
,
.CAHBLTllOI
(
HTRANS_M0
)
,
.CAHBLTO0OI
(
HWRITE_M0
)
,
.CAHBLTII
(
REMAP_M0
)
,
.CAHBLTI0OI
(
HRESP_M0
)
,
.CAHBLTl0OI
(
HRDATA_M0
)
,
.CAHBLTO1OI
(
CAHBLTI1Oll
)
,
.CAHBLTI1OI
(
{
CAHBLTO0IOI
,
CAHBLTl1OOI
,
CAHBLTIIOOI
,
CAHBLTO011
,
CAHBLTl101
,
CAHBLTII01
,
CAHBLTO0l1
,
CAHBLTl1I1
,
CAHBLTIII1
,
CAHBLTO0O1
,
CAHBLTl110
,
CAHBLTII10
,
CAHBLTO000
,
CAHBLTl1l0
,
CAHBLTIIl0
,
CAHBLTO0I0
,
CAHBLTl1O0
}
)
,
.CAHBLTl1OI
(
{
CAHBLTI0IOI
,
CAHBLTOOIOI
,
CAHBLTlIOOI
,
CAHBLTI011
,
CAHBLTOO11
,
CAHBLTlI01
,
CAHBLTI0l1
,
CAHBLTOOl1
,
CAHBLTlII1
,
CAHBLTI0O1
,
CAHBLTOOO1
,
CAHBLTlI10
,
CAHBLTI000
,
CAHBLTOO00
,
CAHBLTlIl0
,
CAHBLTI0I0
,
CAHBLTOOI0
}
)
,
.CAHBLTOOII
(
{
CAHBLTl0IOI
,
CAHBLTIOIOI
,
CAHBLTOlOOI
,
CAHBLTl011
,
CAHBLTIO11
,
CAHBLTOl01
,
CAHBLTl0l1
,
CAHBLTIOl1
,
CAHBLTOlI1
,
CAHBLTl0O1
,
CAHBLTIOO1
,
CAHBLTOl10
,
CAHBLTl000
,
CAHBLTIO00
,
CAHBLTOll0
,
CAHBLTl0I0
,
CAHBLTIOI0
}
)
,
.CAHBLTIOII
(
CAHBLTI11I
)
,
.CAHBLTlOII
(
CAHBLTlI0
)
,
.CAHBLTOIII
(
CAHBLTl11I
)
,
.CAHBLTIIII
(
CAHBLTOOOl
)
,
.CAHBLTlIII
(
CAHBLTIOOl
)
,
.CAHBLTOlII
(
{
CAHBLTlOIOI
,
CAHBLTIlOOI
,
CAHBLTO111
,
CAHBLTlO11
,
CAHBLTIl01
,
CAHBLTO1l1
,
CAHBLTlOl1
,
CAHBLTIlI1
,
CAHBLTO1O1
,
CAHBLTlOO1
,
CAHBLTIl10
,
CAHBLTO100
,
CAHBLTlO00
,
CAHBLTIll0
,
CAHBLTO1I0
,
CAHBLTlOI0
,
CAHBLTIlO0
}
)
,
.CAHBLTIlII
(
{
CAHBLTOIIOI
,
CAHBLTllOOI
,
CAHBLTI111
,
CAHBLTOI11
,
CAHBLTll01
,
CAHBLTI1l1
,
CAHBLTOIl1
,
CAHBLTllI1
,
CAHBLTI1O1
,
CAHBLTOIO1
,
CAHBLTll10
,
CAHBLTI100
,
CAHBLTOI00
,
CAHBLTlll0
,
CAHBLTI1I0
,
CAHBLTOII0
,
CAHBLTllO0
}
)
,
.CAHBLTllII
(
CAHBLTOlO0
)
,
.HRDATA_S0
(
CAHBLTOI0lI
)
,
.HREADYOUT_S0
(
CAHBLTIlO0I
)
,
.HRDATA_S1
(
CAHBLTII0lI
)
,
.HREADYOUT_S1
(
CAHBLTllO0I
)
,
.HRDATA_S2
(
CAHBLTlI0lI
)
,
.HREADYOUT_S2
(
CAHBLTO0O0I
)
,
.HRDATA_S3
(
CAHBLTOl0lI
)
,
.HREADYOUT_S3
(
CAHBLTI0O0I
)
,
.HRDATA_S4
(
CAHBLTIl0lI
)
,
.HREADYOUT_S4
(
CAHBLTl0O0I
)
,
.HRDATA_S5
(
CAHBLTll0lI
)
,
.HREADYOUT_S5
(
CAHBLTO1O0I
)
,
.HRDATA_S6
(
CAHBLTO00lI
)
,
.HREADYOUT_S6
(
CAHBLTI1O0I
)
,
.HRDATA_S7
(
CAHBLTI00lI
)
,
.HREADYOUT_S7
(
CAHBLTl1O0I
)
,
.HRDATA_S8
(
CAHBLTl00lI
)
,
.HREADYOUT_S8
(
CAHBLTOOI0I
)
,
.HRDATA_S9
(
CAHBLTO10lI
)
,
.HREADYOUT_S9
(
CAHBLTIOI0I
)
,
.HRDATA_S10
(
CAHBLTI10lI
)
,
.HREADYOUT_S10
(
CAHBLTlOI0I
)
,
.HRDATA_S11
(
CAHBLTl10lI
)
,
.HREADYOUT_S11
(
CAHBLTOII0I
)
,
.HRDATA_S12
(
CAHBLTOO1lI
)
,
.HREADYOUT_S12
(
CAHBLTIII0I
)
,
.HRDATA_S13
(
CAHBLTIO1lI
)
,
.HREADYOUT_S13
(
CAHBLTlII0I
)
,
.HRDATA_S14
(
CAHBLTlO1lI
)
,
.HREADYOUT_S14
(
CAHBLTOlI0I
)
,
.HRDATA_S15
(
CAHBLTOI1lI
)
,
.HREADYOUT_S15
(
CAHBLTIlI0I
)
,
.HRDATA_S16
(
CAHBLTII1lI
)
,
.HREADYOUT_S16
(
CAHBLTllI0I
)
)
;
CAHBLTIIOI
#
(
.MEMSPACE
(
MEMSPACE
)
,
.HADDR_SHG_CFG
(
HADDR_SHG_CFG
)
,
.CAHBLTI
(
CAHBLTI
)
,
.CAHBLTl
(
CAHBLTlIO0
)
,
.SYNC_RESET
(
SYNC_RESET
)
)
CAHBLTIOIll
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.CAHBLTII
(
1
'b
0
)
,
.CAHBLTlIOI
(
HADDR_M1
)
,
.CAHBLTOlOI
(
HMASTLOCK_M1
)
,
.CAHBLTIlOI
(
HSIZE_M1
)
,
.CAHBLTllOI
(
HTRANS_M1
)
,
.CAHBLTO0OI
(
HWRITE_M1
)
,
.CAHBLTI0OI
(
HRESP_M1
)
,
.CAHBLTl0OI
(
HRDATA_M1
)
,
.CAHBLTO1OI
(
CAHBLTl1Oll
)
,
.CAHBLTI1OI
(
{
CAHBLTOO0lI
,
CAHBLTlIllI
,
CAHBLTI0IlI
,
CAHBLTOOIlI
,
CAHBLTlIOlI
,
CAHBLTI01II
,
CAHBLTOO1II
,
CAHBLTlI0II
,
CAHBLTI0lII
,
CAHBLTOOlII
,
CAHBLTlIIII
,
CAHBLTI0OII
,
CAHBLTOOOII
,
CAHBLTlI1OI
,
CAHBLTI00OI
,
CAHBLTOO0OI
,
CAHBLTlIlOI
}
)
,
.CAHBLTl1OI
(
{
CAHBLTIO0lI
,
CAHBLTOlllI
,
CAHBLTl0IlI
,
CAHBLTIOIlI
,
CAHBLTOlOlI
,
CAHBLTl01II
,
CAHBLTIO1II
,
CAHBLTOl0II
,
CAHBLTl0lII
,
CAHBLTIOlII
,
CAHBLTOlIII
,
CAHBLTl0OII
,
CAHBLTIOOII
,
CAHBLTOl1OI
,
CAHBLTl00OI
,
CAHBLTIO0OI
,
CAHBLTOllOI
}
)
,
.CAHBLTOOII
(
{
CAHBLTlO0lI
,
CAHBLTIlllI
,
CAHBLTO1IlI
,
CAHBLTlOIlI
,
CAHBLTIlOlI
,
CAHBLTO11II
,
CAHBLTlO1II
,
CAHBLTIl0II
,
CAHBLTO1lII
,
CAHBLTlOlII
,
CAHBLTIlIII
,
CAHBLTO1OII
,
CAHBLTlOOII
,
CAHBLTIl1OI
,
CAHBLTO10OI
,
CAHBLTlO0OI
,
CAHBLTIllOI
}
)
,
.CAHBLTIOII
(
CAHBLTlOOl
)
,
.CAHBLTlOII
(
CAHBLTOl0
)
,
.CAHBLTOIII
(
CAHBLTOIOl
)
,
.CAHBLTIIII
(
CAHBLTIIOl
)
,
.CAHBLTlIII
(
CAHBLTlIOl
)
,
.CAHBLTOlII
(
{
CAHBLTllllI
,
CAHBLTI1IlI
,
CAHBLTOIIlI
,
CAHBLTllOlI
,
CAHBLTI11II
,
CAHBLTOI1II
,
CAHBLTll0II
,
CAHBLTI1lII
,
CAHBLTOIlII
,
CAHBLTllIII
,
CAHBLTI1OII
,
CAHBLTOIOII
,
CAHBLTll1OI
,
CAHBLTI10OI
,
CAHBLTOI0OI
,
CAHBLTlllOI
,
CAHBLTI1IOI
}
)
,
.CAHBLTIlII
(
{
CAHBLTO0llI
,
CAHBLTl1IlI
,
CAHBLTIIIlI
,
CAHBLTO0OlI
,
CAHBLTl11II
,
CAHBLTII1II
,
CAHBLTO00II
,
CAHBLTl1lII
,
CAHBLTIIlII
,
CAHBLTO0III
,
CAHBLTl1OII
,
CAHBLTIIOII
,
CAHBLTO01OI
,
CAHBLTl10OI
,
CAHBLTII0OI
,
CAHBLTO0lOI
,
CAHBLTl1IOI
}
)
,
.CAHBLTllII
(
CAHBLTO1IOI
)
,
.HRDATA_S0
(
CAHBLTlI1lI
)
,
.HREADYOUT_S0
(
CAHBLTO0I0I
)
,
.HRDATA_S1
(
CAHBLTOl1lI
)
,
.HREADYOUT_S1
(
CAHBLTI0I0I
)
,
.HRDATA_S2
(
CAHBLTIl1lI
)
,
.HREADYOUT_S2
(
CAHBLTl0I0I
)
,
.HRDATA_S3
(
CAHBLTll1lI
)
,
.HREADYOUT_S3
(
CAHBLTO1I0I
)
,
.HRDATA_S4
(
CAHBLTO01lI
)
,
.HREADYOUT_S4
(
CAHBLTI1I0I
)
,
.HRDATA_S5
(
CAHBLTI01lI
)
,
.HREADYOUT_S5
(
CAHBLTl1I0I
)
,
.HRDATA_S6
(
CAHBLTl01lI
)
,
.HREADYOUT_S6
(
CAHBLTOOl0I
)
,
.HRDATA_S7
(
CAHBLTO11lI
)
,
.HREADYOUT_S7
(
CAHBLTIOl0I
)
,
.HRDATA_S8
(
CAHBLTI11lI
)
,
.HREADYOUT_S8
(
CAHBLTlOl0I
)
,
.HRDATA_S9
(
CAHBLTl11lI
)
,
.HREADYOUT_S9
(
CAHBLTOIl0I
)
,
.HRDATA_S10
(
CAHBLTOOO0I
)
,
.HREADYOUT_S10
(
CAHBLTIIl0I
)
,
.HRDATA_S11
(
CAHBLTIOO0I
)
,
.HREADYOUT_S11
(
CAHBLTlIl0I
)
,
.HRDATA_S12
(
CAHBLTlOO0I
)
,
.HREADYOUT_S12
(
CAHBLTOll0I
)
,
.HRDATA_S13
(
CAHBLTOIO0I
)
,
.HREADYOUT_S13
(
CAHBLTIll0I
)
,
.HRDATA_S14
(
CAHBLTIIO0I
)
,
.HREADYOUT_S14
(
CAHBLTlll0I
)
,
.HRDATA_S15
(
CAHBLTlIO0I
)
,
.HREADYOUT_S15
(
CAHBLTO0l0I
)
,
.HRDATA_S16
(
CAHBLTOlO0I
)
,
.HREADYOUT_S16
(
CAHBLTI0l0I
)
)
;
CAHBLTIIOI
#
(
.MEMSPACE
(
MEMSPACE
)
,
.HADDR_SHG_CFG
(
HADDR_SHG_CFG
)
,
.CAHBLTI
(
CAHBLTI
)
,
.CAHBLTl
(
CAHBLTlIlll
)
,
.SYNC_RESET
(
SYNC_RESET
)
)
CAHBLTO1OI1
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.CAHBLTII
(
1
'b
0
)
,
.CAHBLTlIOI
(
HADDR_M2
)
,
.CAHBLTOlOI
(
HMASTLOCK_M2
)
,
.CAHBLTIlOI
(
HSIZE_M2
)
,
.CAHBLTllOI
(
HTRANS_M2
)
,
.CAHBLTO0OI
(
HWRITE_M2
)
,
.CAHBLTI0OI
(
HRESP_M2
)
,
.CAHBLTl0OI
(
HRDATA_M2
)
,
.CAHBLTO1OI
(
CAHBLTI0OI1
)
,
.CAHBLTI1OI
(
{
CAHBLTI001l
,
CAHBLTOO01l
,
CAHBLTlIl1l
,
CAHBLTI0I1l
,
CAHBLTOOI1l
,
CAHBLTlIO1l
,
CAHBLTI010l
,
CAHBLTOO10l
,
CAHBLTlI00l
,
CAHBLTI0l0l
,
CAHBLTOOl0l
,
CAHBLTlII0l
,
CAHBLTI0O0l
,
CAHBLTOOO0l
,
CAHBLTlI1ll
,
CAHBLTI00ll
,
CAHBLTOO0ll
}
)
,
.CAHBLTl1OI
(
{
CAHBLTl001l
,
CAHBLTIO01l
,
CAHBLTOll1l
,
CAHBLTl0I1l
,
CAHBLTIOI1l
,
CAHBLTOlO1l
,
CAHBLTl010l
,
CAHBLTIO10l
,
CAHBLTOl00l
,
CAHBLTl0l0l
,
CAHBLTIOl0l
,
CAHBLTOlI0l
,
CAHBLTl0O0l
,
CAHBLTIOO0l
,
CAHBLTOl1ll
,
CAHBLTl00ll
,
CAHBLTIO0ll
}
)
,
.CAHBLTOOII
(
{
CAHBLTO101l
,
CAHBLTlO01l
,
CAHBLTIll1l
,
CAHBLTO1I1l
,
CAHBLTlOI1l
,
CAHBLTIlO1l
,
CAHBLTO110l
,
CAHBLTlO10l
,
CAHBLTIl00l
,
CAHBLTO1l0l
,
CAHBLTlOl0l
,
CAHBLTIlI0l
,
CAHBLTO1O0l
,
CAHBLTlOO0l
,
CAHBLTIl1ll
,
CAHBLTO10ll
,
CAHBLTlO0ll
}
)
,
.CAHBLTIOII
(
CAHBLTOlOl
)
,
.CAHBLTlOII
(
CAHBLTIl0
)
,
.CAHBLTOIII
(
CAHBLTIlOl
)
,
.CAHBLTIIII
(
CAHBLTllOl
)
,
.CAHBLTlIII
(
CAHBLTO0Ol
)
,
.CAHBLTOlII
(
{
CAHBLTOI01l
,
CAHBLTlll1l
,
CAHBLTI1I1l
,
CAHBLTOII1l
,
CAHBLTllO1l
,
CAHBLTI110l
,
CAHBLTOI10l
,
CAHBLTll00l
,
CAHBLTI1l0l
,
CAHBLTOIl0l
,
CAHBLTllI0l
,
CAHBLTI1O0l
,
CAHBLTOIO0l
,
CAHBLTll1ll
,
CAHBLTI10ll
,
CAHBLTOI0ll
,
CAHBLTlllll
}
)
,
.CAHBLTIlII
(
{
CAHBLTII01l
,
CAHBLTO0l1l
,
CAHBLTl1I1l
,
CAHBLTIII1l
,
CAHBLTO0O1l
,
CAHBLTl110l
,
CAHBLTII10l
,
CAHBLTO000l
,
CAHBLTl1l0l
,
CAHBLTIIl0l
,
CAHBLTO0I0l
,
CAHBLTl1O0l
,
CAHBLTIIO0l
,
CAHBLTO01ll
,
CAHBLTl10ll
,
CAHBLTII0ll
,
CAHBLTO0lll
}
)
,
.CAHBLTllII
(
CAHBLTIllll
)
,
.HRDATA_S0
(
CAHBLTIIOl0
)
,
.HREADYOUT_S0
(
CAHBLTllll0
)
,
.HRDATA_S1
(
CAHBLTlIOl0
)
,
.HREADYOUT_S1
(
CAHBLTO0ll0
)
,
.HRDATA_S2
(
CAHBLTOlOl0
)
,
.HREADYOUT_S2
(
CAHBLTI0ll0
)
,
.HRDATA_S3
(
CAHBLTIlOl0
)
,
.HREADYOUT_S3
(
CAHBLTl0ll0
)
,
.HRDATA_S4
(
CAHBLTllOl0
)
,
.HREADYOUT_S4
(
CAHBLTO1ll0
)
,
.HRDATA_S5
(
CAHBLTO0Ol0
)
,
.HREADYOUT_S5
(
CAHBLTI1ll0
)
,
.HRDATA_S6
(
CAHBLTI0Ol0
)
,
.HREADYOUT_S6
(
CAHBLTl1ll0
)
,
.HRDATA_S7
(
CAHBLTl0Ol0
)
,
.HREADYOUT_S7
(
CAHBLTOO0l0
)
,
.HRDATA_S8
(
CAHBLTO1Ol0
)
,
.HREADYOUT_S8
(
CAHBLTIO0l0
)
,
.HRDATA_S9
(
CAHBLTI1Ol0
)
,
.HREADYOUT_S9
(
CAHBLTlO0l0
)
,
.HRDATA_S10
(
CAHBLTl1Ol0
)
,
.HREADYOUT_S10
(
CAHBLTOI0l0
)
,
.HRDATA_S11
(
CAHBLTOOIl0
)
,
.HREADYOUT_S11
(
CAHBLTII0l0
)
,
.HRDATA_S12
(
CAHBLTIOIl0
)
,
.HREADYOUT_S12
(
CAHBLTlI0l0
)
,
.HRDATA_S13
(
CAHBLTlOIl0
)
,
.HREADYOUT_S13
(
CAHBLTOl0l0
)
,
.HRDATA_S14
(
CAHBLTOIIl0
)
,
.HREADYOUT_S14
(
CAHBLTIl0l0
)
,
.HRDATA_S15
(
CAHBLTIIIl0
)
,
.HREADYOUT_S15
(
CAHBLTll0l0
)
,
.HRDATA_S16
(
CAHBLTlIIl0
)
,
.HREADYOUT_S16
(
CAHBLTO00l0
)
)
;
CAHBLTIIOI
#
(
.MEMSPACE
(
MEMSPACE
)
,
.HADDR_SHG_CFG
(
HADDR_SHG_CFG
)
,
.CAHBLTI
(
CAHBLTI
)
,
.CAHBLTl
(
CAHBLTOllll
)
,
.SYNC_RESET
(
SYNC_RESET
)
)
CAHBLTI1OI1
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.CAHBLTII
(
1
'b
0
)
,
.CAHBLTlIOI
(
HADDR_M3
)
,
.CAHBLTOlOI
(
HMASTLOCK_M3
)
,
.CAHBLTIlOI
(
HSIZE_M3
)
,
.CAHBLTllOI
(
HTRANS_M3
)
,
.CAHBLTO0OI
(
HWRITE_M3
)
,
.CAHBLTI0OI
(
HRESP_M3
)
,
.CAHBLTl0OI
(
HRDATA_M3
)
,
.CAHBLTO1OI
(
CAHBLTl0OI1
)
,
.CAHBLTI1OI
(
{
CAHBLTIOOl0
,
CAHBLTOl1I0
,
CAHBLTl00I0
,
CAHBLTIO0I0
,
CAHBLTOllI0
,
CAHBLTl0II0
,
CAHBLTIOII0
,
CAHBLTOlOI0
,
CAHBLTl01O0
,
CAHBLTIO1O0
,
CAHBLTOl0O0
,
CAHBLTl0lO0
,
CAHBLTIOlO0
,
CAHBLTOlIO0
,
CAHBLTl0OO0
,
CAHBLTIOOO0
,
CAHBLTOl11l
}
)
,
.CAHBLTl1OI
(
{
CAHBLTlOOl0
,
CAHBLTIl1I0
,
CAHBLTO10I0
,
CAHBLTlO0I0
,
CAHBLTIllI0
,
CAHBLTO1II0
,
CAHBLTlOII0
,
CAHBLTIlOI0
,
CAHBLTO11O0
,
CAHBLTlO1O0
,
CAHBLTIl0O0
,
CAHBLTO1lO0
,
CAHBLTlOlO0
,
CAHBLTIlIO0
,
CAHBLTO1OO0
,
CAHBLTlOOO0
,
CAHBLTIl11l
}
)
,
.CAHBLTOOII
(
{
CAHBLTOIOl0
,
CAHBLTll1I0
,
CAHBLTI10I0
,
CAHBLTOI0I0
,
CAHBLTlllI0
,
CAHBLTI1II0
,
CAHBLTOIII0
,
CAHBLTllOI0
,
CAHBLTI11O0
,
CAHBLTOI1O0
,
CAHBLTll0O0
,
CAHBLTI1lO0
,
CAHBLTOIlO0
,
CAHBLTllIO0
,
CAHBLTI1OO0
,
CAHBLTOIOO0
,
CAHBLTll11l
}
)
,
.CAHBLTIOII
(
CAHBLTI0Ol
)
,
.CAHBLTlOII
(
CAHBLTll0
)
,
.CAHBLTOIII
(
CAHBLTl0Ol
)
,
.CAHBLTIIII
(
CAHBLTO1Ol
)
,
.CAHBLTlIII
(
CAHBLTI1Ol
)
,
.CAHBLTOlII
(
{
CAHBLTO01I0
,
CAHBLTl10I0
,
CAHBLTII0I0
,
CAHBLTO0lI0
,
CAHBLTl1II0
,
CAHBLTIIII0
,
CAHBLTO0OI0
,
CAHBLTl11O0
,
CAHBLTII1O0
,
CAHBLTO00O0
,
CAHBLTl1lO0
,
CAHBLTIIlO0
,
CAHBLTO0IO0
,
CAHBLTl1OO0
,
CAHBLTIIOO0
,
CAHBLTO011l
,
CAHBLTl101l
}
)
,
.CAHBLTIlII
(
{
CAHBLTI01I0
,
CAHBLTOO1I0
,
CAHBLTlI0I0
,
CAHBLTI0lI0
,
CAHBLTOOlI0
,
CAHBLTlIII0
,
CAHBLTI0OI0
,
CAHBLTOOOI0
,
CAHBLTlI1O0
,
CAHBLTI00O0
,
CAHBLTOO0O0
,
CAHBLTlIlO0
,
CAHBLTI0IO0
,
CAHBLTOOIO0
,
CAHBLTlIOO0
,
CAHBLTI011l
,
CAHBLTOO11l
}
)
,
.CAHBLTllII
(
CAHBLTI101l
)
,
.HRDATA_S0
(
CAHBLTOlIl0
)
,
.HREADYOUT_S0
(
CAHBLTI00l0
)
,
.HRDATA_S1
(
CAHBLTIlIl0
)
,
.HREADYOUT_S1
(
CAHBLTl00l0
)
,
.HRDATA_S2
(
CAHBLTllIl0
)
,
.HREADYOUT_S2
(
CAHBLTO10l0
)
,
.HRDATA_S3
(
CAHBLTO0Il0
)
,
.HREADYOUT_S3
(
CAHBLTI10l0
)
,
.HRDATA_S4
(
CAHBLTI0Il0
)
,
.HREADYOUT_S4
(
CAHBLTl10l0
)
,
.HRDATA_S5
(
CAHBLTl0Il0
)
,
.HREADYOUT_S5
(
CAHBLTOO1l0
)
,
.HRDATA_S6
(
CAHBLTO1Il0
)
,
.HREADYOUT_S6
(
CAHBLTIO1l0
)
,
.HRDATA_S7
(
CAHBLTI1Il0
)
,
.HREADYOUT_S7
(
CAHBLTlO1l0
)
,
.HRDATA_S8
(
CAHBLTl1Il0
)
,
.HREADYOUT_S8
(
CAHBLTOI1l0
)
,
.HRDATA_S9
(
CAHBLTOOll0
)
,
.HREADYOUT_S9
(
CAHBLTII1l0
)
,
.HRDATA_S10
(
CAHBLTIOll0
)
,
.HREADYOUT_S10
(
CAHBLTlI1l0
)
,
.HRDATA_S11
(
CAHBLTlOll0
)
,
.HREADYOUT_S11
(
CAHBLTOl1l0
)
,
.HRDATA_S12
(
CAHBLTOIll0
)
,
.HREADYOUT_S12
(
CAHBLTIl1l0
)
,
.HRDATA_S13
(
CAHBLTIIll0
)
,
.HREADYOUT_S13
(
CAHBLTll1l0
)
,
.HRDATA_S14
(
CAHBLTlIll0
)
,
.HREADYOUT_S14
(
CAHBLTO01l0
)
,
.HRDATA_S15
(
CAHBLTOlll0
)
,
.HREADYOUT_S15
(
CAHBLTI01l0
)
,
.HRDATA_S16
(
CAHBLTIlll0
)
,
.HREADYOUT_S16
(
CAHBLTl01l0
)
)
;
CAHBLTOI1I
#
(
.SYNC_RESET
(
SYNC_RESET
)
)
CAHBLTlOIll
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.CAHBLTII1I
(
CAHBLTl0l0I
)
,
.CAHBLTI0OI
(
CAHBLTI100I
)
,
.CAHBLTlI1I
(
HSEL_S0
)
,
.CAHBLTlIOI
(
HADDR_S0
)
,
.CAHBLTIlOI
(
HSIZE_S0
)
,
.CAHBLTllOI
(
HTRANS_S0
)
,
.CAHBLTO0OI
(
HWRITE_S0
)
,
.CAHBLTOl1I
(
HWDATA_S0
)
,
.CAHBLTIl1I
(
HREADY_S0
)
,
.CAHBLTOlOI
(
HMASTLOCK_S0
)
,
.CAHBLTOI0
(
{
CAHBLTII11l
,
CAHBLTI1lll
,
CAHBLTOIlOI
,
CAHBLTO1O0
}
)
,
.CAHBLTll1I
(
{
CAHBLTlI11l
,
CAHBLTl1lll
,
CAHBLTIIlOI
,
CAHBLTI1O0
}
)
,
.CAHBLTO01I
(
{
CAHBLTll1O1
,
CAHBLTOl0O1
,
CAHBLTl01Il
,
CAHBLTO00Il
}
)
,
.CAHBLTI01I
(
{
CAHBLTIO11l
,
CAHBLTI0lll
,
CAHBLTOOlOI
,
CAHBLTO0O0
}
)
,
.CAHBLTl01I
(
{
CAHBLTlO11l
,
CAHBLTl0lll
,
CAHBLTIOlOI
,
CAHBLTI0O0
}
)
,
.CAHBLTO11I
(
{
CAHBLTOI11l
,
CAHBLTO1lll
,
CAHBLTlOlOI
,
CAHBLTl0O0
}
)
,
.CAHBLTI11I
(
CAHBLTIIl1I
)
,
.CAHBLTlI0
(
CAHBLTO1IOl
)
,
.CAHBLTl11I
(
CAHBLTll11I
)
,
.CAHBLTOOOl
(
CAHBLTIO1Ol
)
,
.CAHBLTIOOl
(
CAHBLTlIIIl
)
,
.CAHBLTlOOl
(
CAHBLTOl01I
)
,
.CAHBLTOl0
(
CAHBLTl1lOl
)
,
.CAHBLTOIOl
(
CAHBLTI0OOl
)
,
.CAHBLTIIOl
(
CAHBLTOIOIl
)
,
.CAHBLTlIOl
(
CAHBLTIllIl
)
,
.CAHBLTOlOl
(
CAHBLTIOl00
)
,
.CAHBLTIl0
(
CAHBLTO0I10
)
,
.CAHBLTIlOl
(
CAHBLTlI100
)
,
.CAHBLTllOl
(
CAHBLTI1010
)
,
.CAHBLTO0Ol
(
CAHBLTlOIO1
)
,
.CAHBLTI0Ol
(
CAHBLTOI000
)
,
.CAHBLTll0
(
CAHBLTl0l10
)
,
.CAHBLTl0Ol
(
CAHBLTIlO10
)
,
.CAHBLTO1Ol
(
CAHBLTOOOO1
)
,
.CAHBLTI1Ol
(
CAHBLTIIlO1
)
,
.HWDATA_M0
(
CAHBLTOOO1I
)
,
.HWDATA_M1
(
CAHBLTlOI1I
)
,
.HWDATA_M2
(
CAHBLTO11l0
)
,
.HWDATA_M3
(
CAHBLTl1O00
)
)
;
CAHBLTOI1I
#
(
.SYNC_RESET
(
SYNC_RESET
)
)
CAHBLTOIIll
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.CAHBLTII1I
(
CAHBLTO1l0I
)
,
.CAHBLTI0OI
(
CAHBLTl100I
)
,
.CAHBLTlI1I
(
HSEL_S1
)
,
.CAHBLTlIOI
(
HADDR_S1
)
,
.CAHBLTIlOI
(
HSIZE_S1
)
,
.CAHBLTllOI
(
HTRANS_S1
)
,
.CAHBLTO0OI
(
HWRITE_S1
)
,
.CAHBLTOl1I
(
HWDATA_S1
)
,
.CAHBLTIl1I
(
HREADY_S1
)
,
.CAHBLTOlOI
(
HMASTLOCK_S1
)
,
.CAHBLTOI0
(
{
CAHBLTl111l
,
CAHBLTll0ll
,
CAHBLTI1lOI
,
CAHBLTIlI0
}
)
,
.CAHBLTll1I
(
{
CAHBLTOOOO0
,
CAHBLTO00ll
,
CAHBLTl1lOI
,
CAHBLTllI0
}
)
,
.CAHBLTO01I
(
{
CAHBLTO01O1
,
CAHBLTIl0O1
,
CAHBLTO11Il
,
CAHBLTI00Il
}
)
,
.CAHBLTI01I
(
{
CAHBLTl011l
,
CAHBLTlI0ll
,
CAHBLTI0lOI
,
CAHBLTIII0
}
)
,
.CAHBLTl01I
(
{
CAHBLTO111l
,
CAHBLTOl0ll
,
CAHBLTl0lOI
,
CAHBLTlII0
}
)
,
.CAHBLTO11I
(
{
CAHBLTI111l
,
CAHBLTIl0ll
,
CAHBLTO1lOI
,
CAHBLTOlI0
}
)
,
.CAHBLTI11I
(
CAHBLTlIl1I
)
,
.CAHBLTlI0
(
CAHBLTI1IOl
)
,
.CAHBLTl11I
(
CAHBLTO011I
)
,
.CAHBLTOOOl
(
CAHBLTlO1Ol
)
,
.CAHBLTIOOl
(
CAHBLTOlIIl
)
,
.CAHBLTlOOl
(
CAHBLTIl01I
)
,
.CAHBLTOl0
(
CAHBLTOO0Ol
)
,
.CAHBLTOIOl
(
CAHBLTl0OOl
)
,
.CAHBLTIIOl
(
CAHBLTIIOIl
)
,
.CAHBLTlIOl
(
CAHBLTlllIl
)
,
.CAHBLTOlOl
(
CAHBLTlOl00
)
,
.CAHBLTIl0
(
CAHBLTI0I10
)
,
.CAHBLTIlOl
(
CAHBLTOl100
)
,
.CAHBLTllOl
(
CAHBLTl1010
)
,
.CAHBLTO0Ol
(
CAHBLTOIIO1
)
,
.CAHBLTI0Ol
(
CAHBLTII000
)
,
.CAHBLTll0
(
CAHBLTO1l10
)
,
.CAHBLTl0Ol
(
CAHBLTllO10
)
,
.CAHBLTO1Ol
(
CAHBLTIOOO1
)
,
.CAHBLTI1Ol
(
CAHBLTlIlO1
)
,
.HWDATA_M0
(
CAHBLTIOO1I
)
,
.HWDATA_M1
(
CAHBLTOII1I
)
,
.HWDATA_M2
(
CAHBLTI11l0
)
,
.HWDATA_M3
(
CAHBLTOOI00
)
)
;
CAHBLTOI1I
#
(
.SYNC_RESET
(
SYNC_RESET
)
)
CAHBLTIIIll
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.CAHBLTII1I
(
CAHBLTI1l0I
)
,
.CAHBLTI0OI
(
CAHBLTOO10I
)
,
.CAHBLTlI1I
(
HSEL_S2
)
,
.CAHBLTlIOI
(
HADDR_S2
)
,
.CAHBLTIlOI
(
HSIZE_S2
)
,
.CAHBLTllOI
(
HTRANS_S2
)
,
.CAHBLTO0OI
(
HWRITE_S2
)
,
.CAHBLTOl1I
(
HWDATA_S2
)
,
.CAHBLTIl1I
(
HREADY_S2
)
,
.CAHBLTOlOI
(
HMASTLOCK_S2
)
,
.CAHBLTOI0
(
{
CAHBLTO0OO0
,
CAHBLTOI1ll
,
CAHBLTll0OI
,
CAHBLTlOl0
}
)
,
.CAHBLTll1I
(
{
CAHBLTI0OO0
,
CAHBLTII1ll
,
CAHBLTO00OI
,
CAHBLTOIl0
}
)
,
.CAHBLTO01I
(
{
CAHBLTI01O1
,
CAHBLTll0O1
,
CAHBLTI11Il
,
CAHBLTl00Il
}
)
,
.CAHBLTI01I
(
{
CAHBLTOlOO0
,
CAHBLTOO1ll
,
CAHBLTlI0OI
,
CAHBLTl1I0
}
)
,
.CAHBLTl01I
(
{
CAHBLTIlOO0
,
CAHBLTIO1ll
,
CAHBLTOl0OI
,
CAHBLTOOl0
}
)
,
.CAHBLTO11I
(
{
CAHBLTllOO0
,
CAHBLTlO1ll
,
CAHBLTIl0OI
,
CAHBLTIOl0
}
)
,
.CAHBLTI11I
(
CAHBLTOll1I
)
,
.CAHBLTlI0
(
CAHBLTl1IOl
)
,
.CAHBLTl11I
(
CAHBLTI011I
)
,
.CAHBLTOOOl
(
CAHBLTOI1Ol
)
,
.CAHBLTIOOl
(
CAHBLTIlIIl
)
,
.CAHBLTlOOl
(
CAHBLTll01I
)
,
.CAHBLTOl0
(
CAHBLTIO0Ol
)
,
.CAHBLTOIOl
(
CAHBLTO1OOl
)
,
.CAHBLTIIOl
(
CAHBLTlIOIl
)
,
.CAHBLTlIOl
(
CAHBLTO0lIl
)
,
.CAHBLTOlOl
(
CAHBLTOIl00
)
,
.CAHBLTIl0
(
CAHBLTl0I10
)
,
.CAHBLTIlOl
(
CAHBLTIl100
)
,
.CAHBLTllOl
(
CAHBLTOO110
)
,
.CAHBLTO0Ol
(
CAHBLTIIIO1
)
,
.CAHBLTI0Ol
(
CAHBLTlI000
)
,
.CAHBLTll0
(
CAHBLTI1l10
)
,
.CAHBLTl0Ol
(
CAHBLTO0O10
)
,
.CAHBLTO1Ol
(
CAHBLTlOOO1
)
,
.CAHBLTI1Ol
(
CAHBLTOllO1
)
,
.HWDATA_M0
(
CAHBLTlOO1I
)
,
.HWDATA_M1
(
CAHBLTIII1I
)
,
.HWDATA_M2
(
CAHBLTl11l0
)
,
.HWDATA_M3
(
CAHBLTIOI00
)
)
;
CAHBLTOI1I
#
(
.SYNC_RESET
(
SYNC_RESET
)
)
CAHBLTlIIll
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.CAHBLTII1I
(
CAHBLTl1l0I
)
,
.CAHBLTI0OI
(
CAHBLTIO10I
)
,
.CAHBLTlI1I
(
HSEL_S3
)
,
.CAHBLTlIOI
(
HADDR_S3
)
,
.CAHBLTIlOI
(
HSIZE_S3
)
,
.CAHBLTllOI
(
HTRANS_S3
)
,
.CAHBLTO0OI
(
HWRITE_S3
)
,
.CAHBLTOl1I
(
HWDATA_S3
)
,
.CAHBLTIl1I
(
HREADY_S3
)
,
.CAHBLTOlOI
(
HMASTLOCK_S3
)
,
.CAHBLTOI0
(
{
CAHBLTIIIO0
,
CAHBLTI11ll
,
CAHBLTOI1OI
,
CAHBLTO1l0
}
)
,
.CAHBLTll1I
(
{
CAHBLTlIIO0
,
CAHBLTl11ll
,
CAHBLTII1OI
,
CAHBLTI1l0
}
)
,
.CAHBLTO01I
(
{
CAHBLTl01O1
,
CAHBLTO00O1
,
CAHBLTl11Il
,
CAHBLTO10Il
}
)
,
.CAHBLTI01I
(
{
CAHBLTIOIO0
,
CAHBLTI01ll
,
CAHBLTOO1OI
,
CAHBLTO0l0
}
)
,
.CAHBLTl01I
(
{
CAHBLTlOIO0
,
CAHBLTl01ll
,
CAHBLTIO1OI
,
CAHBLTI0l0
}
)
,
.CAHBLTO11I
(
{
CAHBLTOIIO0
,
CAHBLTO11ll
,
CAHBLTlO1OI
,
CAHBLTl0l0
}
)
,
.CAHBLTI11I
(
CAHBLTIll1I
)
,
.CAHBLTlI0
(
CAHBLTOOlOl
)
,
.CAHBLTl11I
(
CAHBLTl011I
)
,
.CAHBLTOOOl
(
CAHBLTII1Ol
)
,
.CAHBLTIOOl
(
CAHBLTllIIl
)
,
.CAHBLTlOOl
(
CAHBLTO001I
)
,
.CAHBLTOl0
(
CAHBLTlO0Ol
)
,
.CAHBLTOIOl
(
CAHBLTI1OOl
)
,
.CAHBLTIIOl
(
CAHBLTOlOIl
)
,
.CAHBLTlIOl
(
CAHBLTI0lIl
)
,
.CAHBLTOlOl
(
CAHBLTIIl00
)
,
.CAHBLTIl0
(
CAHBLTO1I10
)
,
.CAHBLTIlOl
(
CAHBLTll100
)
,
.CAHBLTllOl
(
CAHBLTIO110
)
,
.CAHBLTO0Ol
(
CAHBLTlIIO1
)
,
.CAHBLTI0Ol
(
CAHBLTOl000
)
,
.CAHBLTll0
(
CAHBLTl1l10
)
,
.CAHBLTl0Ol
(
CAHBLTI0O10
)
,
.CAHBLTO1Ol
(
CAHBLTOIOO1
)
,
.CAHBLTI1Ol
(
CAHBLTIllO1
)
,
.HWDATA_M0
(
CAHBLTOIO1I
)
,
.HWDATA_M1
(
CAHBLTlII1I
)
,
.HWDATA_M2
(
CAHBLTOOO00
)
,
.HWDATA_M3
(
CAHBLTlOI00
)
)
;
CAHBLTOI1I
#
(
.SYNC_RESET
(
SYNC_RESET
)
)
CAHBLTOlIll
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.CAHBLTII1I
(
CAHBLTOO00I
)
,
.CAHBLTI0OI
(
CAHBLTlO10I
)
,
.CAHBLTlI1I
(
HSEL_S4
)
,
.CAHBLTlIOI
(
HADDR_S4
)
,
.CAHBLTIlOI
(
HSIZE_S4
)
,
.CAHBLTllOI
(
HTRANS_S4
)
,
.CAHBLTO0OI
(
HWRITE_S4
)
,
.CAHBLTOl1I
(
HWDATA_S4
)
,
.CAHBLTIl1I
(
HREADY_S4
)
,
.CAHBLTOlOI
(
HMASTLOCK_S4
)
,
.CAHBLTOI0
(
{
CAHBLTl1IO0
,
CAHBLTllO0l
,
CAHBLTI11OI
,
CAHBLTIl00
}
)
,
.CAHBLTll1I
(
{
CAHBLTOOlO0
,
CAHBLTO0O0l
,
CAHBLTl11OI
,
CAHBLTll00
}
)
,
.CAHBLTO01I
(
{
CAHBLTO11O1
,
CAHBLTI00O1
,
CAHBLTOOOll
,
CAHBLTI10Il
}
)
,
.CAHBLTI01I
(
{
CAHBLTl0IO0
,
CAHBLTlIO0l
,
CAHBLTI01OI
,
CAHBLTII00
}
)
,
.CAHBLTl01I
(
{
CAHBLTO1IO0
,
CAHBLTOlO0l
,
CAHBLTl01OI
,
CAHBLTlI00
}
)
,
.CAHBLTO11I
(
{
CAHBLTI1IO0
,
CAHBLTIlO0l
,
CAHBLTO11OI
,
CAHBLTOl00
}
)
,
.CAHBLTI11I
(
CAHBLTlll1I
)
,
.CAHBLTlI0
(
CAHBLTIOlOl
)
,
.CAHBLTl11I
(
CAHBLTO111I
)
,
.CAHBLTOOOl
(
CAHBLTlI1Ol
)
,
.CAHBLTIOOl
(
CAHBLTO0IIl
)
,
.CAHBLTlOOl
(
CAHBLTI001I
)
,
.CAHBLTOl0
(
CAHBLTOI0Ol
)
,
.CAHBLTOIOl
(
CAHBLTl1OOl
)
,
.CAHBLTIIOl
(
CAHBLTIlOIl
)
,
.CAHBLTlIOl
(
CAHBLTl0lIl
)
,
.CAHBLTOlOl
(
CAHBLTlIl00
)
,
.CAHBLTIl0
(
CAHBLTI1I10
)
,
.CAHBLTIlOl
(
CAHBLTO0100
)
,
.CAHBLTllOl
(
CAHBLTlO110
)
,
.CAHBLTO0Ol
(
CAHBLTOlIO1
)
,
.CAHBLTI0Ol
(
CAHBLTIl000
)
,
.CAHBLTll0
(
CAHBLTOO010
)
,
.CAHBLTl0Ol
(
CAHBLTl0O10
)
,
.CAHBLTO1Ol
(
CAHBLTIIOO1
)
,
.CAHBLTI1Ol
(
CAHBLTlllO1
)
,
.HWDATA_M0
(
CAHBLTIIO1I
)
,
.HWDATA_M1
(
CAHBLTOlI1I
)
,
.HWDATA_M2
(
CAHBLTIOO00
)
,
.HWDATA_M3
(
CAHBLTOII00
)
)
;
CAHBLTOI1I
#
(
.SYNC_RESET
(
SYNC_RESET
)
)
CAHBLTIlIll
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.CAHBLTII1I
(
CAHBLTIO00I
)
,
.CAHBLTI0OI
(
CAHBLTOI10I
)
,
.CAHBLTlI1I
(
HSEL_S5
)
,
.CAHBLTlIOI
(
HADDR_S5
)
,
.CAHBLTIlOI
(
HSIZE_S5
)
,
.CAHBLTllOI
(
HTRANS_S5
)
,
.CAHBLTO0OI
(
HWRITE_S5
)
,
.CAHBLTOl1I
(
HWDATA_S5
)
,
.CAHBLTIl1I
(
HREADY_S5
)
,
.CAHBLTOlOI
(
HMASTLOCK_S5
)
,
.CAHBLTOI0
(
{
CAHBLTO0lO0
,
CAHBLTOII0l
,
CAHBLTllOII
,
CAHBLTlO10
}
)
,
.CAHBLTll1I
(
{
CAHBLTI0lO0
,
CAHBLTIII0l
,
CAHBLTO0OII
,
CAHBLTOI10
}
)
,
.CAHBLTO01I
(
{
CAHBLTI11O1
,
CAHBLTl00O1
,
CAHBLTIOOll
,
CAHBLTl10Il
}
)
,
.CAHBLTI01I
(
{
CAHBLTOllO0
,
CAHBLTOOI0l
,
CAHBLTlIOII
,
CAHBLTl100
}
)
,
.CAHBLTl01I
(
{
CAHBLTIllO0
,
CAHBLTIOI0l
,
CAHBLTOlOII
,
CAHBLTOO10
}
)
,
.CAHBLTO11I
(
{
CAHBLTlllO0
,
CAHBLTlOI0l
,
CAHBLTIlOII
,
CAHBLTIO10
}
)
,
.CAHBLTI11I
(
CAHBLTO0l1I
)
,
.CAHBLTlI0
(
CAHBLTlOlOl
)
,
.CAHBLTl11I
(
CAHBLTI111I
)
,
.CAHBLTOOOl
(
CAHBLTOl1Ol
)
,
.CAHBLTIOOl
(
CAHBLTI0IIl
)
,
.CAHBLTlOOl
(
CAHBLTl001I
)
,
.CAHBLTOl0
(
CAHBLTII0Ol
)
,
.CAHBLTOIOl
(
CAHBLTOOIOl
)
,
.CAHBLTIIOl
(
CAHBLTllOIl
)
,
.CAHBLTlIOl
(
CAHBLTO1lIl
)
,
.CAHBLTOlOl
(
CAHBLTOll00
)
,
.CAHBLTIl0
(
CAHBLTl1I10
)
,
.CAHBLTIlOl
(
CAHBLTI0100
)
,
.CAHBLTllOl
(
CAHBLTOI110
)
,
.CAHBLTO0Ol
(
CAHBLTIlIO1
)
,
.CAHBLTI0Ol
(
CAHBLTll000
)
,
.CAHBLTll0
(
CAHBLTIO010
)
,
.CAHBLTl0Ol
(
CAHBLTO1O10
)
,
.CAHBLTO1Ol
(
CAHBLTlIOO1
)
,
.CAHBLTI1Ol
(
CAHBLTO0lO1
)
,
.HWDATA_M0
(
CAHBLTlIO1I
)
,
.HWDATA_M1
(
CAHBLTIlI1I
)
,
.HWDATA_M2
(
CAHBLTlOO00
)
,
.HWDATA_M3
(
CAHBLTIII00
)
)
;
CAHBLTOI1I
#
(
.SYNC_RESET
(
SYNC_RESET
)
)
CAHBLTllIll
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.CAHBLTII1I
(
CAHBLTlO00I
)
,
.CAHBLTI0OI
(
CAHBLTII10I
)
,
.CAHBLTlI1I
(
HSEL_S6
)
,
.CAHBLTlIOI
(
HADDR_S6
)
,
.CAHBLTIlOI
(
HSIZE_S6
)
,
.CAHBLTllOI
(
HTRANS_S6
)
,
.CAHBLTO0OI
(
HWRITE_S6
)
,
.CAHBLTOl1I
(
HWDATA_S6
)
,
.CAHBLTIl1I
(
HREADY_S6
)
,
.CAHBLTOlOI
(
HMASTLOCK_S6
)
,
.CAHBLTOI0
(
{
CAHBLTII0O0
,
CAHBLTI1I0l
,
CAHBLTOIIII
,
CAHBLTO110
}
)
,
.CAHBLTll1I
(
{
CAHBLTlI0O0
,
CAHBLTl1I0l
,
CAHBLTIIIII
,
CAHBLTI110
}
)
,
.CAHBLTO01I
(
{
CAHBLTl11O1
,
CAHBLTO10O1
,
CAHBLTlOOll
,
CAHBLTOO1Il
}
)
,
.CAHBLTI01I
(
{
CAHBLTIO0O0
,
CAHBLTI0I0l
,
CAHBLTOOIII
,
CAHBLTO010
}
)
,
.CAHBLTl01I
(
{
CAHBLTlO0O0
,
CAHBLTl0I0l
,
CAHBLTIOIII
,
CAHBLTI010
}
)
,
.CAHBLTO11I
(
{
CAHBLTOI0O0
,
CAHBLTO1I0l
,
CAHBLTlOIII
,
CAHBLTl010
}
)
,
.CAHBLTI11I
(
CAHBLTI0l1I
)
,
.CAHBLTlI0
(
CAHBLTOIlOl
)
,
.CAHBLTl11I
(
CAHBLTl111I
)
,
.CAHBLTOOOl
(
CAHBLTIl1Ol
)
,
.CAHBLTIOOl
(
CAHBLTl0IIl
)
,
.CAHBLTlOOl
(
CAHBLTO101I
)
,
.CAHBLTOl0
(
CAHBLTlI0Ol
)
,
.CAHBLTOIOl
(
CAHBLTIOIOl
)
,
.CAHBLTIIOl
(
CAHBLTO0OIl
)
,
.CAHBLTlIOl
(
CAHBLTI1lIl
)
,
.CAHBLTOlOl
(
CAHBLTIll00
)
,
.CAHBLTIl0
(
CAHBLTOOl10
)
,
.CAHBLTIlOl
(
CAHBLTl0100
)
,
.CAHBLTllOl
(
CAHBLTII110
)
,
.CAHBLTO0Ol
(
CAHBLTllIO1
)
,
.CAHBLTI0Ol
(
CAHBLTO0000
)
,
.CAHBLTll0
(
CAHBLTlO010
)
,
.CAHBLTl0Ol
(
CAHBLTI1O10
)
,
.CAHBLTO1Ol
(
CAHBLTOlOO1
)
,
.CAHBLTI1Ol
(
CAHBLTI0lO1
)
,
.HWDATA_M0
(
CAHBLTOlO1I
)
,
.HWDATA_M1
(
CAHBLTllI1I
)
,
.HWDATA_M2
(
CAHBLTOIO00
)
,
.HWDATA_M3
(
CAHBLTlII00
)
)
;
CAHBLTOI1I
#
(
.SYNC_RESET
(
SYNC_RESET
)
)
CAHBLTO0Ill
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.CAHBLTII1I
(
CAHBLTOI00I
)
,
.CAHBLTI0OI
(
CAHBLTlI10I
)
,
.CAHBLTlI1I
(
HSEL_S7
)
,
.CAHBLTlIOI
(
HADDR_S7
)
,
.CAHBLTIlOI
(
HSIZE_S7
)
,
.CAHBLTllOI
(
HTRANS_S7
)
,
.CAHBLTO0OI
(
HWRITE_S7
)
,
.CAHBLTOl1I
(
HWDATA_S7
)
,
.CAHBLTIl1I
(
HREADY_S7
)
,
.CAHBLTOlOI
(
HMASTLOCK_S7
)
,
.CAHBLTOI0
(
{
CAHBLTl10O0
,
CAHBLTlll0l
,
CAHBLTI1III
,
CAHBLTIlO1
}
)
,
.CAHBLTll1I
(
{
CAHBLTOO1O0
,
CAHBLTO0l0l
,
CAHBLTl1III
,
CAHBLTllO1
}
)
,
.CAHBLTO01I
(
{
CAHBLTOOOI1
,
CAHBLTI10O1
,
CAHBLTOIOll
,
CAHBLTIO1Il
}
)
,
.CAHBLTI01I
(
{
CAHBLTl00O0
,
CAHBLTlIl0l
,
CAHBLTI0III
,
CAHBLTIIO1
}
)
,
.CAHBLTl01I
(
{
CAHBLTO10O0
,
CAHBLTOll0l
,
CAHBLTl0III
,
CAHBLTlIO1
}
)
,
.CAHBLTO11I
(
{
CAHBLTI10O0
,
CAHBLTIll0l
,
CAHBLTO1III
,
CAHBLTOlO1
}
)
,
.CAHBLTI11I
(
CAHBLTl0l1I
)
,
.CAHBLTlI0
(
CAHBLTIIlOl
)
,
.CAHBLTl11I
(
CAHBLTOOOOl
)
,
.CAHBLTOOOl
(
CAHBLTll1Ol
)
,
.CAHBLTIOOl
(
CAHBLTO1IIl
)
,
.CAHBLTlOOl
(
CAHBLTI101I
)
,
.CAHBLTOl0
(
CAHBLTOl0Ol
)
,
.CAHBLTOIOl
(
CAHBLTlOIOl
)
,
.CAHBLTIIOl
(
CAHBLTI0OIl
)
,
.CAHBLTlIOl
(
CAHBLTl1lIl
)
,
.CAHBLTOlOl
(
CAHBLTlll00
)
,
.CAHBLTIl0
(
CAHBLTIOl10
)
,
.CAHBLTIlOl
(
CAHBLTO1100
)
,
.CAHBLTllOl
(
CAHBLTlI110
)
,
.CAHBLTO0Ol
(
CAHBLTO0IO1
)
,
.CAHBLTI0Ol
(
CAHBLTI0000
)
,
.CAHBLTll0
(
CAHBLTOI010
)
,
.CAHBLTl0Ol
(
CAHBLTl1O10
)
,
.CAHBLTO1Ol
(
CAHBLTIlOO1
)
,
.CAHBLTI1Ol
(
CAHBLTl0lO1
)
,
.HWDATA_M0
(
CAHBLTIlO1I
)
,
.HWDATA_M1
(
CAHBLTO0I1I
)
,
.HWDATA_M2
(
CAHBLTIIO00
)
,
.HWDATA_M3
(
CAHBLTOlI00
)
)
;
CAHBLTOI1I
#
(
.SYNC_RESET
(
SYNC_RESET
)
)
CAHBLTI0Ill
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.CAHBLTII1I
(
CAHBLTII00I
)
,
.CAHBLTI0OI
(
CAHBLTOl10I
)
,
.CAHBLTlI1I
(
HSEL_S8
)
,
.CAHBLTlIOI
(
HADDR_S8
)
,
.CAHBLTIlOI
(
HSIZE_S8
)
,
.CAHBLTllOI
(
HTRANS_S8
)
,
.CAHBLTO0OI
(
HWRITE_S8
)
,
.CAHBLTOl1I
(
HWDATA_S8
)
,
.CAHBLTIl1I
(
HREADY_S8
)
,
.CAHBLTOlOI
(
HMASTLOCK_S8
)
,
.CAHBLTOI0
(
{
CAHBLTO01O0
,
CAHBLTOI00l
,
CAHBLTlllII
,
CAHBLTlOI1
}
)
,
.CAHBLTll1I
(
{
CAHBLTI01O0
,
CAHBLTII00l
,
CAHBLTO0lII
,
CAHBLTOII1
}
)
,
.CAHBLTO01I
(
{
CAHBLTIOOI1
,
CAHBLTl10O1
,
CAHBLTIIOll
,
CAHBLTlO1Il
}
)
,
.CAHBLTI01I
(
{
CAHBLTOl1O0
,
CAHBLTOO00l
,
CAHBLTlIlII
,
CAHBLTl1O1
}
)
,
.CAHBLTl01I
(
{
CAHBLTIl1O0
,
CAHBLTIO00l
,
CAHBLTOllII
,
CAHBLTOOI1
}
)
,
.CAHBLTO11I
(
{
CAHBLTll1O0
,
CAHBLTlO00l
,
CAHBLTIllII
,
CAHBLTIOI1
}
)
,
.CAHBLTI11I
(
CAHBLTO1l1I
)
,
.CAHBLTlI0
(
CAHBLTlIlOl
)
,
.CAHBLTl11I
(
CAHBLTIOOOl
)
,
.CAHBLTOOOl
(
CAHBLTO01Ol
)
,
.CAHBLTIOOl
(
CAHBLTI1IIl
)
,
.CAHBLTlOOl
(
CAHBLTl101I
)
,
.CAHBLTOl0
(
CAHBLTIl0Ol
)
,
.CAHBLTOIOl
(
CAHBLTOIIOl
)
,
.CAHBLTIIOl
(
CAHBLTl0OIl
)
,
.CAHBLTlIOl
(
CAHBLTOO0Il
)
,
.CAHBLTOlOl
(
CAHBLTO0l00
)
,
.CAHBLTIl0
(
CAHBLTlOl10
)
,
.CAHBLTIlOl
(
CAHBLTI1100
)
,
.CAHBLTllOl
(
CAHBLTOl110
)
,
.CAHBLTO0Ol
(
CAHBLTI0IO1
)
,
.CAHBLTI0Ol
(
CAHBLTl0000
)
,
.CAHBLTll0
(
CAHBLTII010
)
,
.CAHBLTl0Ol
(
CAHBLTOOI10
)
,
.CAHBLTO1Ol
(
CAHBLTllOO1
)
,
.CAHBLTI1Ol
(
CAHBLTO1lO1
)
,
.HWDATA_M0
(
CAHBLTllO1I
)
,
.HWDATA_M1
(
CAHBLTI0I1I
)
,
.HWDATA_M2
(
CAHBLTlIO00
)
,
.HWDATA_M3
(
CAHBLTIlI00
)
)
;
CAHBLTOI1I
#
(
.SYNC_RESET
(
SYNC_RESET
)
)
CAHBLTl0Ill
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.CAHBLTII1I
(
CAHBLTlI00I
)
,
.CAHBLTI0OI
(
CAHBLTIl10I
)
,
.CAHBLTlI1I
(
HSEL_S9
)
,
.CAHBLTlIOI
(
HADDR_S9
)
,
.CAHBLTIlOI
(
HSIZE_S9
)
,
.CAHBLTllOI
(
HTRANS_S9
)
,
.CAHBLTO0OI
(
HWRITE_S9
)
,
.CAHBLTOl1I
(
HWDATA_S9
)
,
.CAHBLTIl1I
(
HREADY_S9
)
,
.CAHBLTOlOI
(
HMASTLOCK_S9
)
,
.CAHBLTOI0
(
{
CAHBLTIIOI0
,
CAHBLTI100l
,
CAHBLTOI0II
,
CAHBLTO1I1
}
)
,
.CAHBLTll1I
(
{
CAHBLTlIOI0
,
CAHBLTl100l
,
CAHBLTII0II
,
CAHBLTI1I1
}
)
,
.CAHBLTO01I
(
{
CAHBLTlOOI1
,
CAHBLTOO1O1
,
CAHBLTlIOll
,
CAHBLTOI1Il
}
)
,
.CAHBLTI01I
(
{
CAHBLTIOOI0
,
CAHBLTI000l
,
CAHBLTOO0II
,
CAHBLTO0I1
}
)
,
.CAHBLTl01I
(
{
CAHBLTlOOI0
,
CAHBLTl000l
,
CAHBLTIO0II
,
CAHBLTI0I1
}
)
,
.CAHBLTO11I
(
{
CAHBLTOIOI0
,
CAHBLTO100l
,
CAHBLTlO0II
,
CAHBLTl0I1
}
)
,
.CAHBLTI11I
(
CAHBLTI1l1I
)
,
.CAHBLTlI0
(
CAHBLTOllOl
)
,
.CAHBLTl11I
(
CAHBLTlOOOl
)
,
.CAHBLTOOOl
(
CAHBLTI01Ol
)
,
.CAHBLTIOOl
(
CAHBLTl1IIl
)
,
.CAHBLTlOOl
(
CAHBLTOO11I
)
,
.CAHBLTOl0
(
CAHBLTll0Ol
)
,
.CAHBLTOIOl
(
CAHBLTIIIOl
)
,
.CAHBLTIIOl
(
CAHBLTO1OIl
)
,
.CAHBLTlIOl
(
CAHBLTIO0Il
)
,
.CAHBLTOlOl
(
CAHBLTI0l00
)
,
.CAHBLTIl0
(
CAHBLTOIl10
)
,
.CAHBLTIlOl
(
CAHBLTl1100
)
,
.CAHBLTllOl
(
CAHBLTIl110
)
,
.CAHBLTO0Ol
(
CAHBLTl0IO1
)
,
.CAHBLTI0Ol
(
CAHBLTO1000
)
,
.CAHBLTll0
(
CAHBLTlI010
)
,
.CAHBLTl0Ol
(
CAHBLTIOI10
)
,
.CAHBLTO1Ol
(
CAHBLTO0OO1
)
,
.CAHBLTI1Ol
(
CAHBLTI1lO1
)
,
.HWDATA_M0
(
CAHBLTO0O1I
)
,
.HWDATA_M1
(
CAHBLTl0I1I
)
,
.HWDATA_M2
(
CAHBLTOlO00
)
,
.HWDATA_M3
(
CAHBLTllI00
)
)
;
CAHBLTOI1I
#
(
.SYNC_RESET
(
SYNC_RESET
)
)
CAHBLTO1Ill
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.CAHBLTII1I
(
CAHBLTOl00I
)
,
.CAHBLTI0OI
(
CAHBLTll10I
)
,
.CAHBLTlI1I
(
HSEL_S10
)
,
.CAHBLTlIOI
(
HADDR_S10
)
,
.CAHBLTIlOI
(
HSIZE_S10
)
,
.CAHBLTllOI
(
HTRANS_S10
)
,
.CAHBLTO0OI
(
HWRITE_S10
)
,
.CAHBLTOl1I
(
HWDATA_S10
)
,
.CAHBLTIl1I
(
HREADY_S10
)
,
.CAHBLTOlOI
(
HMASTLOCK_S10
)
,
.CAHBLTOI0
(
{
CAHBLTl1OI0
,
CAHBLTll10l
,
CAHBLTI10II
,
CAHBLTIll1
}
)
,
.CAHBLTll1I
(
{
CAHBLTOOII0
,
CAHBLTO010l
,
CAHBLTl10II
,
CAHBLTlll1
}
)
,
.CAHBLTO01I
(
{
CAHBLTOIOI1
,
CAHBLTIO1O1
,
CAHBLTOlOll
,
CAHBLTII1Il
}
)
,
.CAHBLTI01I
(
{
CAHBLTl0OI0
,
CAHBLTlI10l
,
CAHBLTI00II
,
CAHBLTIIl1
}
)
,
.CAHBLTl01I
(
{
CAHBLTO1OI0
,
CAHBLTOl10l
,
CAHBLTl00II
,
CAHBLTlIl1
}
)
,
.CAHBLTO11I
(
{
CAHBLTI1OI0
,
CAHBLTIl10l
,
CAHBLTO10II
,
CAHBLTOll1
}
)
,
.CAHBLTI11I
(
CAHBLTl1l1I
)
,
.CAHBLTlI0
(
CAHBLTIllOl
)
,
.CAHBLTl11I
(
CAHBLTOIOOl
)
,
.CAHBLTOOOl
(
CAHBLTl01Ol
)
,
.CAHBLTIOOl
(
CAHBLTOOlIl
)
,
.CAHBLTlOOl
(
CAHBLTIO11I
)
,
.CAHBLTOl0
(
CAHBLTO00Ol
)
,
.CAHBLTOIOl
(
CAHBLTlIIOl
)
,
.CAHBLTIIOl
(
CAHBLTI1OIl
)
,
.CAHBLTlIOl
(
CAHBLTlO0Il
)
,
.CAHBLTOlOl
(
CAHBLTl0l00
)
,
.CAHBLTIl0
(
CAHBLTIIl10
)
,
.CAHBLTIlOl
(
CAHBLTOOO10
)
,
.CAHBLTllOl
(
CAHBLTll110
)
,
.CAHBLTO0Ol
(
CAHBLTO1IO1
)
,
.CAHBLTI0Ol
(
CAHBLTI1000
)
,
.CAHBLTll0
(
CAHBLTOl010
)
,
.CAHBLTl0Ol
(
CAHBLTlOI10
)
,
.CAHBLTO1Ol
(
CAHBLTI0OO1
)
,
.CAHBLTI1Ol
(
CAHBLTl1lO1
)
,
.HWDATA_M0
(
CAHBLTI0O1I
)
,
.HWDATA_M1
(
CAHBLTO1I1I
)
,
.HWDATA_M2
(
CAHBLTIlO00
)
,
.HWDATA_M3
(
CAHBLTO0I00
)
)
;
CAHBLTOI1I
#
(
.SYNC_RESET
(
SYNC_RESET
)
)
CAHBLTI1Ill
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.CAHBLTII1I
(
CAHBLTIl00I
)
,
.CAHBLTI0OI
(
CAHBLTO010I
)
,
.CAHBLTlI1I
(
HSEL_S11
)
,
.CAHBLTlIOI
(
HADDR_S11
)
,
.CAHBLTIlOI
(
HSIZE_S11
)
,
.CAHBLTllOI
(
HTRANS_S11
)
,
.CAHBLTO0OI
(
HWRITE_S11
)
,
.CAHBLTOl1I
(
HWDATA_S11
)
,
.CAHBLTIl1I
(
HREADY_S11
)
,
.CAHBLTOlOI
(
HMASTLOCK_S11
)
,
.CAHBLTOI0
(
{
CAHBLTO0II0
,
CAHBLTOIO1l
,
CAHBLTll1II
,
CAHBLTlO01
}
)
,
.CAHBLTll1I
(
{
CAHBLTI0II0
,
CAHBLTIIO1l
,
CAHBLTO01II
,
CAHBLTOI01
}
)
,
.CAHBLTO01I
(
{
CAHBLTIIOI1
,
CAHBLTlO1O1
,
CAHBLTIlOll
,
CAHBLTlI1Il
}
)
,
.CAHBLTI01I
(
{
CAHBLTOlII0
,
CAHBLTOOO1l
,
CAHBLTlI1II
,
CAHBLTl1l1
}
)
,
.CAHBLTl01I
(
{
CAHBLTIlII0
,
CAHBLTIOO1l
,
CAHBLTOl1II
,
CAHBLTOO01
}
)
,
.CAHBLTO11I
(
{
CAHBLTllII0
,
CAHBLTlOO1l
,
CAHBLTIl1II
,
CAHBLTIO01
}
)
,
.CAHBLTI11I
(
CAHBLTOO01I
)
,
.CAHBLTlI0
(
CAHBLTlllOl
)
,
.CAHBLTl11I
(
CAHBLTIIOOl
)
,
.CAHBLTOOOl
(
CAHBLTO11Ol
)
,
.CAHBLTIOOl
(
CAHBLTIOlIl
)
,
.CAHBLTlOOl
(
CAHBLTlO11I
)
,
.CAHBLTOl0
(
CAHBLTI00Ol
)
,
.CAHBLTOIOl
(
CAHBLTOlIOl
)
,
.CAHBLTIIOl
(
CAHBLTl1OIl
)
,
.CAHBLTlIOl
(
CAHBLTOI0Il
)
,
.CAHBLTOlOl
(
CAHBLTO1l00
)
,
.CAHBLTIl0
(
CAHBLTlIl10
)
,
.CAHBLTIlOl
(
CAHBLTIOO10
)
,
.CAHBLTllOl
(
CAHBLTO0110
)
,
.CAHBLTO0Ol
(
CAHBLTI1IO1
)
,
.CAHBLTI0Ol
(
CAHBLTl1000
)
,
.CAHBLTll0
(
CAHBLTIl010
)
,
.CAHBLTl0Ol
(
CAHBLTOII10
)
,
.CAHBLTO1Ol
(
CAHBLTl0OO1
)
,
.CAHBLTI1Ol
(
CAHBLTOO0O1
)
,
.HWDATA_M0
(
CAHBLTl0O1I
)
,
.HWDATA_M1
(
CAHBLTI1I1I
)
,
.HWDATA_M2
(
CAHBLTllO00
)
,
.HWDATA_M3
(
CAHBLTI0I00
)
)
;
CAHBLTOI1I
#
(
.SYNC_RESET
(
SYNC_RESET
)
)
CAHBLTl1Ill
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.CAHBLTII1I
(
CAHBLTll00I
)
,
.CAHBLTI0OI
(
CAHBLTI010I
)
,
.CAHBLTlI1I
(
HSEL_S12
)
,
.CAHBLTlIOI
(
HADDR_S12
)
,
.CAHBLTIlOI
(
HSIZE_S12
)
,
.CAHBLTllOI
(
HTRANS_S12
)
,
.CAHBLTO0OI
(
HWRITE_S12
)
,
.CAHBLTOl1I
(
HWDATA_S12
)
,
.CAHBLTIl1I
(
HREADY_S12
)
,
.CAHBLTOlOI
(
HMASTLOCK_S12
)
,
.CAHBLTOI0
(
{
CAHBLTIIlI0
,
CAHBLTI1O1l
,
CAHBLTOIOlI
,
CAHBLTO101
}
)
,
.CAHBLTll1I
(
{
CAHBLTlIlI0
,
CAHBLTl1O1l
,
CAHBLTIIOlI
,
CAHBLTI101
}
)
,
.CAHBLTO01I
(
{
CAHBLTlIOI1
,
CAHBLTOI1O1
,
CAHBLTllOll
,
CAHBLTOl1Il
}
)
,
.CAHBLTI01I
(
{
CAHBLTIOlI0
,
CAHBLTI0O1l
,
CAHBLTOOOlI
,
CAHBLTO001
}
)
,
.CAHBLTl01I
(
{
CAHBLTlOlI0
,
CAHBLTl0O1l
,
CAHBLTIOOlI
,
CAHBLTI001
}
)
,
.CAHBLTO11I
(
{
CAHBLTOIlI0
,
CAHBLTO1O1l
,
CAHBLTlOOlI
,
CAHBLTl001
}
)
,
.CAHBLTI11I
(
CAHBLTIO01I
)
,
.CAHBLTlI0
(
CAHBLTO0lOl
)
,
.CAHBLTl11I
(
CAHBLTlIOOl
)
,
.CAHBLTOOOl
(
CAHBLTI11Ol
)
,
.CAHBLTIOOl
(
CAHBLTlOlIl
)
,
.CAHBLTlOOl
(
CAHBLTOI11I
)
,
.CAHBLTOl0
(
CAHBLTl00Ol
)
,
.CAHBLTOIOl
(
CAHBLTIlIOl
)
,
.CAHBLTIIOl
(
CAHBLTOOIIl
)
,
.CAHBLTlIOl
(
CAHBLTII0Il
)
,
.CAHBLTOlOl
(
CAHBLTI1l00
)
,
.CAHBLTIl0
(
CAHBLTOll10
)
,
.CAHBLTIlOl
(
CAHBLTlOO10
)
,
.CAHBLTllOl
(
CAHBLTI0110
)
,
.CAHBLTO0Ol
(
CAHBLTl1IO1
)
,
.CAHBLTI0Ol
(
CAHBLTOO100
)
,
.CAHBLTll0
(
CAHBLTll010
)
,
.CAHBLTl0Ol
(
CAHBLTIII10
)
,
.CAHBLTO1Ol
(
CAHBLTO1OO1
)
,
.CAHBLTI1Ol
(
CAHBLTIO0O1
)
,
.HWDATA_M0
(
CAHBLTO1O1I
)
,
.HWDATA_M1
(
CAHBLTl1I1I
)
,
.HWDATA_M2
(
CAHBLTO0O00
)
,
.HWDATA_M3
(
CAHBLTl0I00
)
)
;
CAHBLTOI1I
#
(
.SYNC_RESET
(
SYNC_RESET
)
)
CAHBLTOOlll
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.CAHBLTII1I
(
CAHBLTO000I
)
,
.CAHBLTI0OI
(
CAHBLTl010I
)
,
.CAHBLTlI1I
(
HSEL_S13
)
,
.CAHBLTlIOI
(
HADDR_S13
)
,
.CAHBLTIlOI
(
HSIZE_S13
)
,
.CAHBLTllOI
(
HTRANS_S13
)
,
.CAHBLTO0OI
(
HWRITE_S13
)
,
.CAHBLTOl1I
(
HWDATA_S13
)
,
.CAHBLTIl1I
(
HREADY_S13
)
,
.CAHBLTOlOI
(
HMASTLOCK_S13
)
,
.CAHBLTOI0
(
{
CAHBLTl1lI0
,
CAHBLTllI1l
,
CAHBLTI1OlI
,
CAHBLTIl11
}
)
,
.CAHBLTll1I
(
{
CAHBLTOO0I0
,
CAHBLTO0I1l
,
CAHBLTl1OlI
,
CAHBLTll11
}
)
,
.CAHBLTO01I
(
{
CAHBLTOlOI1
,
CAHBLTII1O1
,
CAHBLTO0Oll
,
CAHBLTIl1Il
}
)
,
.CAHBLTI01I
(
{
CAHBLTl0lI0
,
CAHBLTlII1l
,
CAHBLTI0OlI
,
CAHBLTII11
}
)
,
.CAHBLTl01I
(
{
CAHBLTO1lI0
,
CAHBLTOlI1l
,
CAHBLTl0OlI
,
CAHBLTlI11
}
)
,
.CAHBLTO11I
(
{
CAHBLTI1lI0
,
CAHBLTIlI1l
,
CAHBLTO1OlI
,
CAHBLTOl11
}
)
,
.CAHBLTI11I
(
CAHBLTlO01I
)
,
.CAHBLTlI0
(
CAHBLTI0lOl
)
,
.CAHBLTl11I
(
CAHBLTOlOOl
)
,
.CAHBLTOOOl
(
CAHBLTl11Ol
)
,
.CAHBLTIOOl
(
CAHBLTOIlIl
)
,
.CAHBLTlOOl
(
CAHBLTII11I
)
,
.CAHBLTOl0
(
CAHBLTO10Ol
)
,
.CAHBLTOIOl
(
CAHBLTllIOl
)
,
.CAHBLTIIOl
(
CAHBLTIOIIl
)
,
.CAHBLTlIOl
(
CAHBLTlI0Il
)
,
.CAHBLTOlOl
(
CAHBLTl1l00
)
,
.CAHBLTIl0
(
CAHBLTIll10
)
,
.CAHBLTIlOl
(
CAHBLTOIO10
)
,
.CAHBLTllOl
(
CAHBLTl0110
)
,
.CAHBLTO0Ol
(
CAHBLTOOlO1
)
,
.CAHBLTI0Ol
(
CAHBLTIO100
)
,
.CAHBLTll0
(
CAHBLTO0010
)
,
.CAHBLTl0Ol
(
CAHBLTlII10
)
,
.CAHBLTO1Ol
(
CAHBLTI1OO1
)
,
.CAHBLTI1Ol
(
CAHBLTlO0O1
)
,
.HWDATA_M0
(
CAHBLTI1O1I
)
,
.HWDATA_M1
(
CAHBLTOOl1I
)
,
.HWDATA_M2
(
CAHBLTI0O00
)
,
.HWDATA_M3
(
CAHBLTO1I00
)
)
;
CAHBLTOI1I
#
(
.SYNC_RESET
(
SYNC_RESET
)
)
CAHBLTIOlll
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.CAHBLTII1I
(
CAHBLTI000I
)
,
.CAHBLTI0OI
(
CAHBLTO110I
)
,
.CAHBLTlI1I
(
HSEL_S14
)
,
.CAHBLTlIOI
(
HADDR_S14
)
,
.CAHBLTIlOI
(
HSIZE_S14
)
,
.CAHBLTllOI
(
HTRANS_S14
)
,
.CAHBLTO0OI
(
HWRITE_S14
)
,
.CAHBLTOl1I
(
HWDATA_S14
)
,
.CAHBLTIl1I
(
HREADY_S14
)
,
.CAHBLTOlOI
(
HMASTLOCK_S14
)
,
.CAHBLTOI0
(
{
CAHBLTO00I0
,
CAHBLTOIl1l
,
CAHBLTllIlI
,
CAHBLTlOOOI
}
)
,
.CAHBLTll1I
(
{
CAHBLTI00I0
,
CAHBLTIIl1l
,
CAHBLTO0IlI
,
CAHBLTOIOOI
}
)
,
.CAHBLTO01I
(
{
CAHBLTIlOI1
,
CAHBLTlI1O1
,
CAHBLTI0Oll
,
CAHBLTll1Il
}
)
,
.CAHBLTI01I
(
{
CAHBLTOl0I0
,
CAHBLTOOl1l
,
CAHBLTlIIlI
,
CAHBLTl111
}
)
,
.CAHBLTl01I
(
{
CAHBLTIl0I0
,
CAHBLTIOl1l
,
CAHBLTOlIlI
,
CAHBLTOOOOI
}
)
,
.CAHBLTO11I
(
{
CAHBLTll0I0
,
CAHBLTlOl1l
,
CAHBLTIlIlI
,
CAHBLTIOOOI
}
)
,
.CAHBLTI11I
(
CAHBLTOI01I
)
,
.CAHBLTlI0
(
CAHBLTl0lOl
)
,
.CAHBLTl11I
(
CAHBLTIlOOl
)
,
.CAHBLTOOOl
(
CAHBLTOOOIl
)
,
.CAHBLTIOOl
(
CAHBLTIIlIl
)
,
.CAHBLTlOOl
(
CAHBLTlI11I
)
,
.CAHBLTOl0
(
CAHBLTI10Ol
)
,
.CAHBLTOIOl
(
CAHBLTO0IOl
)
,
.CAHBLTIIOl
(
CAHBLTlOIIl
)
,
.CAHBLTlIOl
(
CAHBLTOl0Il
)
,
.CAHBLTOlOl
(
CAHBLTOO000
)
,
.CAHBLTIl0
(
CAHBLTlll10
)
,
.CAHBLTIlOl
(
CAHBLTIIO10
)
,
.CAHBLTllOl
(
CAHBLTO1110
)
,
.CAHBLTO0Ol
(
CAHBLTIOlO1
)
,
.CAHBLTI0Ol
(
CAHBLTlO100
)
,
.CAHBLTll0
(
CAHBLTI0010
)
,
.CAHBLTl0Ol
(
CAHBLTOlI10
)
,
.CAHBLTO1Ol
(
CAHBLTl1OO1
)
,
.CAHBLTI1Ol
(
CAHBLTOI0O1
)
,
.HWDATA_M0
(
CAHBLTl1O1I
)
,
.HWDATA_M1
(
CAHBLTIOl1I
)
,
.HWDATA_M2
(
CAHBLTl0O00
)
,
.HWDATA_M3
(
CAHBLTI1I00
)
)
;
CAHBLTOI1I
#
(
.SYNC_RESET
(
SYNC_RESET
)
)
CAHBLTlOlll
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.CAHBLTII1I
(
CAHBLTl000I
)
,
.CAHBLTI0OI
(
CAHBLTI110I
)
,
.CAHBLTlI1I
(
HSEL_S15
)
,
.CAHBLTlIOI
(
HADDR_S15
)
,
.CAHBLTIlOI
(
HSIZE_S15
)
,
.CAHBLTllOI
(
HTRANS_S15
)
,
.CAHBLTO0OI
(
HWRITE_S15
)
,
.CAHBLTOl1I
(
HWDATA_S15
)
,
.CAHBLTIl1I
(
HREADY_S15
)
,
.CAHBLTOlOI
(
HMASTLOCK_S15
)
,
.CAHBLTOI0
(
{
CAHBLTII1I0
,
CAHBLTI1l1l
,
CAHBLTOIllI
,
CAHBLTO1OOI
}
)
,
.CAHBLTll1I
(
{
CAHBLTlI1I0
,
CAHBLTl1l1l
,
CAHBLTIIllI
,
CAHBLTI1OOI
}
)
,
.CAHBLTO01I
(
{
CAHBLTllOI1
,
CAHBLTOl1O1
,
CAHBLTl0Oll
,
CAHBLTO01Il
}
)
,
.CAHBLTI01I
(
{
CAHBLTIO1I0
,
CAHBLTI0l1l
,
CAHBLTOOllI
,
CAHBLTO0OOI
}
)
,
.CAHBLTl01I
(
{
CAHBLTlO1I0
,
CAHBLTl0l1l
,
CAHBLTIOllI
,
CAHBLTI0OOI
}
)
,
.CAHBLTO11I
(
{
CAHBLTOI1I0
,
CAHBLTO1l1l
,
CAHBLTlOllI
,
CAHBLTl0OOI
}
)
,
.CAHBLTI11I
(
CAHBLTII01I
)
,
.CAHBLTlI0
(
CAHBLTO1lOl
)
,
.CAHBLTl11I
(
CAHBLTllOOl
)
,
.CAHBLTOOOl
(
CAHBLTIOOIl
)
,
.CAHBLTIOOl
(
CAHBLTlIlIl
)
,
.CAHBLTlOOl
(
CAHBLTOl11I
)
,
.CAHBLTOl0
(
CAHBLTl10Ol
)
,
.CAHBLTOIOl
(
CAHBLTI0IOl
)
,
.CAHBLTIIOl
(
CAHBLTOIIIl
)
,
.CAHBLTlIOl
(
CAHBLTIl0Il
)
,
.CAHBLTOlOl
(
CAHBLTIO000
)
,
.CAHBLTIl0
(
CAHBLTO0l10
)
,
.CAHBLTIlOl
(
CAHBLTlIO10
)
,
.CAHBLTllOl
(
CAHBLTI1110
)
,
.CAHBLTO0Ol
(
CAHBLTlOlO1
)
,
.CAHBLTI0Ol
(
CAHBLTOI100
)
,
.CAHBLTll0
(
CAHBLTl0010
)
,
.CAHBLTl0Ol
(
CAHBLTIlI10
)
,
.CAHBLTO1Ol
(
CAHBLTOOIO1
)
,
.CAHBLTI1Ol
(
CAHBLTII0O1
)
,
.HWDATA_M0
(
CAHBLTOOI1I
)
,
.HWDATA_M1
(
CAHBLTlOl1I
)
,
.HWDATA_M2
(
CAHBLTO1O00
)
,
.HWDATA_M3
(
CAHBLTl1I00
)
)
;
CAHBLTOI1I
#
(
.SYNC_RESET
(
SYNC_RESET
)
)
CAHBLTOIlll
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.CAHBLTII1I
(
CAHBLTO100I
)
,
.CAHBLTI0OI
(
CAHBLTl110I
)
,
.CAHBLTlI1I
(
HSEL_S16
)
,
.CAHBLTlIOI
(
HADDR_S16
)
,
.CAHBLTIlOI
(
HSIZE_S16
)
,
.CAHBLTllOI
(
HTRANS_S16
)
,
.CAHBLTO0OI
(
HWRITE_S16
)
,
.CAHBLTOl1I
(
HWDATA_S16
)
,
.CAHBLTIl1I
(
HREADY_S16
)
,
.CAHBLTOlOI
(
HMASTLOCK_S16
)
,
.CAHBLTOI0
(
{
CAHBLTl11I0
,
CAHBLTll01l
,
CAHBLTI1llI
,
CAHBLTIlIOI
}
)
,
.CAHBLTll1I
(
{
CAHBLTOOOl0
,
CAHBLTO001l
,
CAHBLTl1llI
,
CAHBLTllIOI
}
)
,
.CAHBLTO01I
(
{
CAHBLTO0OI1
,
CAHBLTIl1O1
,
CAHBLTO1Oll
,
CAHBLTI01Il
}
)
,
.CAHBLTI01I
(
{
CAHBLTl01I0
,
CAHBLTlI01l
,
CAHBLTI0llI
,
CAHBLTIIIOI
}
)
,
.CAHBLTl01I
(
{
CAHBLTO11I0
,
CAHBLTOl01l
,
CAHBLTl0llI
,
CAHBLTlIIOI
}
)
,
.CAHBLTO11I
(
{
CAHBLTI11I0
,
CAHBLTIl01l
,
CAHBLTO1llI
,
CAHBLTOlIOI
}
)
,
.CAHBLTI11I
(
CAHBLTlI01I
)
,
.CAHBLTlI0
(
CAHBLTI1lOl
)
,
.CAHBLTl11I
(
CAHBLTO0OOl
)
,
.CAHBLTOOOl
(
CAHBLTlOOIl
)
,
.CAHBLTIOOl
(
CAHBLTOllIl
)
,
.CAHBLTlOOl
(
CAHBLTIl11I
)
,
.CAHBLTOl0
(
CAHBLTOO1Ol
)
,
.CAHBLTOIOl
(
CAHBLTl0IOl
)
,
.CAHBLTIIOl
(
CAHBLTIIIIl
)
,
.CAHBLTlIOl
(
CAHBLTll0Il
)
,
.CAHBLTOlOl
(
CAHBLTlO000
)
,
.CAHBLTIl0
(
CAHBLTI0l10
)
,
.CAHBLTIlOl
(
CAHBLTOlO10
)
,
.CAHBLTllOl
(
CAHBLTl1110
)
,
.CAHBLTO0Ol
(
CAHBLTOIlO1
)
,
.CAHBLTI0Ol
(
CAHBLTII100
)
,
.CAHBLTll0
(
CAHBLTO1010
)
,
.CAHBLTl0Ol
(
CAHBLTllI10
)
,
.CAHBLTO1Ol
(
CAHBLTIOIO1
)
,
.CAHBLTI1Ol
(
CAHBLTlI0O1
)
,
.HWDATA_M0
(
CAHBLTIOI1I
)
,
.HWDATA_M1
(
CAHBLTOIl1I
)
,
.HWDATA_M2
(
CAHBLTI1O00
)
,
.HWDATA_M3
(
CAHBLTOOl00
)
)
;
assign
HREADY_M0
=
CAHBLTI1Oll
;
assign
HREADY_M1
=
CAHBLTl1Oll
;
assign
HREADY_M2
=
CAHBLTI0OI1
;
assign
HREADY_M3
=
CAHBLTl0OI1
;
endmodule
