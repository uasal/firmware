// Actel Corporation Proprietary and Confidential
// Copyright 2013 Actel Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE ACTEL LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
// SVN Revision Information:
// SVN $Revision: 23120 $
// SVN $Date: 2014-07-17 15:26:23 +0100 (Thu, 17 Jul 2014) $
`timescale 1ns/1ps
module
CAHBLTlO0
#
(
parameter
SYNC_RESET
=
0
)
(
input
HCLK,
input
HRESETN,
input
[
3
:
0
]
CAHBLTOI0,
input
CAHBLTII0,
input
CAHBLTlI0,
input
CAHBLTOl0,
input
CAHBLTIl0,
input
CAHBLTll0,
output
reg
[
3
:
0
]
CAHBLTO00
)
;
localparam
CAHBLTI00
=
4
'b
0000
;
localparam
CAHBLTl00
=
4
'b
0001
;
localparam
CAHBLTO10
=
4
'b
0010
;
localparam
CAHBLTI10
=
4
'b
0011
;
localparam
CAHBLTl10
=
4
'b
0100
;
localparam
CAHBLTOO1
=
4
'b
0101
;
localparam
CAHBLTIO1
=
4
'b
0110
;
localparam
CAHBLTlO1
=
4
'b
0111
;
localparam
CAHBLTOI1
=
4
'b
1000
;
localparam
CAHBLTII1
=
4
'b
1001
;
localparam
CAHBLTlI1
=
4
'b
1010
;
localparam
CAHBLTOl1
=
4
'b
1011
;
localparam
CAHBLTIl1
=
4
'b
1100
;
localparam
CAHBLTll1
=
4
'b
1101
;
localparam
CAHBLTO01
=
4
'b
1110
;
localparam
CAHBLTI01
=
4
'b
1111
;
localparam
CAHBLTl01
=
4
'b
0001
;
localparam
CAHBLTO11
=
4
'b
0010
;
localparam
CAHBLTI11
=
4
'b
0100
;
localparam
CAHBLTl11
=
4
'b
1000
;
localparam
CAHBLTOOOI
=
4
'b
0000
;
reg
[
127
:
0
]
CAHBLTIOOI
;
reg
[
3
:
0
]
CAHBLTlOOI
;
reg
[
3
:
0
]
CAHBLTOIOI
;
wire
CAHBLTOO0
;
wire
CAHBLTIO0
;
assign
CAHBLTOO0
=
(
SYNC_RESET
==
1
)
?
1
'b
1
:
HRESETN
;
assign
CAHBLTIO0
=
(
SYNC_RESET
==
1
)
?
HRESETN
:
1
'b
1
;
always
@
(
*
)
begin
CAHBLTO00
=
CAHBLTOOOI
;
case
(
CAHBLTOIOI
)
CAHBLTll1
:
begin
CAHBLTIOOI
=
"M3DONE"
;
if
(
CAHBLTOI0
[
0
]
)
begin
if
(
CAHBLTlI0
)
CAHBLTlOOI
=
CAHBLTO10
;
else
begin
CAHBLTO00
=
CAHBLTl01
;
if
(
CAHBLTII0
)
CAHBLTlOOI
=
CAHBLTl00
;
else
CAHBLTlOOI
=
CAHBLTI00
;
end
end
else
if
(
CAHBLTOI0
[
1
]
)
begin
if
(
CAHBLTOl0
)
CAHBLTlOOI
=
CAHBLTIO1
;
else
begin
CAHBLTO00
=
CAHBLTO11
;
if
(
CAHBLTII0
)
CAHBLTlOOI
=
CAHBLTOO1
;
else
CAHBLTlOOI
=
CAHBLTl10
;
end
end
else
if
(
CAHBLTOI0
[
2
]
)
begin
if
(
CAHBLTIl0
)
CAHBLTlOOI
=
CAHBLTlI1
;
else
begin
CAHBLTO00
=
CAHBLTI11
;
if
(
CAHBLTII0
)
CAHBLTlOOI
=
CAHBLTII1
;
else
CAHBLTlOOI
=
CAHBLTOI1
;
end
end
else
if
(
CAHBLTOI0
[
3
]
)
begin
if
(
CAHBLTll0
)
CAHBLTlOOI
=
CAHBLTO01
;
else
begin
CAHBLTO00
=
CAHBLTl11
;
if
(
CAHBLTII0
)
CAHBLTlOOI
=
CAHBLTll1
;
else
CAHBLTlOOI
=
CAHBLTIl1
;
end
end
else
begin
CAHBLTlOOI
=
CAHBLTll1
;
end
end
CAHBLTII1
:
begin
CAHBLTIOOI
=
"M2DONE"
;
if
(
CAHBLTOI0
[
3
]
)
begin
if
(
CAHBLTll0
)
CAHBLTlOOI
=
CAHBLTO01
;
else
begin
CAHBLTO00
=
CAHBLTl11
;
if
(
CAHBLTII0
)
CAHBLTlOOI
=
CAHBLTll1
;
else
CAHBLTlOOI
=
CAHBLTIl1
;
end
end
else
if
(
CAHBLTOI0
[
0
]
)
begin
if
(
CAHBLTlI0
)
CAHBLTlOOI
=
CAHBLTO10
;
else
begin
CAHBLTO00
=
CAHBLTl01
;
if
(
CAHBLTII0
)
CAHBLTlOOI
=
CAHBLTl00
;
else
CAHBLTlOOI
=
CAHBLTI00
;
end
end
else
if
(
CAHBLTOI0
[
1
]
)
begin
if
(
CAHBLTOl0
)
CAHBLTlOOI
=
CAHBLTIO1
;
else
begin
CAHBLTO00
=
CAHBLTO11
;
if
(
CAHBLTII0
)
CAHBLTlOOI
=
CAHBLTOO1
;
else
CAHBLTlOOI
=
CAHBLTl10
;
end
end
else
if
(
CAHBLTOI0
[
2
]
)
begin
if
(
CAHBLTIl0
)
CAHBLTlOOI
=
CAHBLTlI1
;
else
begin
CAHBLTO00
=
CAHBLTI11
;
if
(
CAHBLTII0
)
CAHBLTlOOI
=
CAHBLTII1
;
else
CAHBLTlOOI
=
CAHBLTOI1
;
end
end
else
begin
CAHBLTlOOI
=
CAHBLTII1
;
end
end
CAHBLTOO1
:
begin
CAHBLTIOOI
=
"M1DONE"
;
if
(
CAHBLTOI0
[
2
]
)
begin
if
(
CAHBLTIl0
)
CAHBLTlOOI
=
CAHBLTlI1
;
else
begin
CAHBLTO00
=
CAHBLTI11
;
if
(
CAHBLTII0
)
CAHBLTlOOI
=
CAHBLTII1
;
else
CAHBLTlOOI
=
CAHBLTOI1
;
end
end
else
if
(
CAHBLTOI0
[
3
]
)
begin
if
(
CAHBLTll0
)
CAHBLTlOOI
=
CAHBLTO01
;
else
begin
CAHBLTO00
=
CAHBLTl11
;
if
(
CAHBLTII0
)
CAHBLTlOOI
=
CAHBLTll1
;
else
CAHBLTlOOI
=
CAHBLTIl1
;
end
end
else
if
(
CAHBLTOI0
[
0
]
)
begin
if
(
CAHBLTlI0
)
CAHBLTlOOI
=
CAHBLTO10
;
else
begin
CAHBLTO00
=
CAHBLTl01
;
if
(
CAHBLTII0
)
CAHBLTlOOI
=
CAHBLTl00
;
else
CAHBLTlOOI
=
CAHBLTI00
;
end
end
else
if
(
CAHBLTOI0
[
1
]
)
begin
if
(
CAHBLTOl0
)
CAHBLTlOOI
=
CAHBLTIO1
;
else
begin
CAHBLTO00
=
CAHBLTO11
;
if
(
CAHBLTII0
)
CAHBLTlOOI
=
CAHBLTOO1
;
else
CAHBLTlOOI
=
CAHBLTl10
;
end
end
else
begin
CAHBLTlOOI
=
CAHBLTOO1
;
end
end
CAHBLTl00
:
begin
CAHBLTIOOI
=
"M0DONE"
;
if
(
CAHBLTOI0
[
1
]
)
begin
if
(
CAHBLTOl0
)
CAHBLTlOOI
=
CAHBLTIO1
;
else
begin
CAHBLTO00
=
CAHBLTO11
;
if
(
CAHBLTII0
)
CAHBLTlOOI
=
CAHBLTOO1
;
else
CAHBLTlOOI
=
CAHBLTl10
;
end
end
else
if
(
CAHBLTOI0
[
2
]
)
begin
if
(
CAHBLTIl0
)
CAHBLTlOOI
=
CAHBLTlI1
;
else
begin
CAHBLTO00
=
CAHBLTI11
;
if
(
CAHBLTII0
)
CAHBLTlOOI
=
CAHBLTII1
;
else
CAHBLTlOOI
=
CAHBLTOI1
;
end
end
else
if
(
CAHBLTOI0
[
3
]
)
begin
if
(
CAHBLTll0
)
CAHBLTlOOI
=
CAHBLTO01
;
else
begin
CAHBLTO00
=
CAHBLTl11
;
if
(
CAHBLTII0
)
CAHBLTlOOI
=
CAHBLTll1
;
else
CAHBLTlOOI
=
CAHBLTIl1
;
end
end
else
if
(
CAHBLTOI0
[
0
]
)
begin
if
(
CAHBLTlI0
)
CAHBLTlOOI
=
CAHBLTO10
;
else
begin
CAHBLTO00
=
CAHBLTl01
;
if
(
CAHBLTII0
)
CAHBLTlOOI
=
CAHBLTl00
;
else
CAHBLTlOOI
=
CAHBLTI00
;
end
end
else
begin
CAHBLTlOOI
=
CAHBLTl00
;
end
end
CAHBLTI00
:
begin
CAHBLTIOOI
=
"M0EXTEND"
;
CAHBLTO00
=
CAHBLTl01
;
if
(
CAHBLTII0
)
CAHBLTlOOI
=
CAHBLTl00
;
else
CAHBLTlOOI
=
CAHBLTI00
;
end
CAHBLTl10
:
begin
CAHBLTIOOI
=
"M1EXTEND"
;
CAHBLTO00
=
CAHBLTO11
;
if
(
CAHBLTII0
)
CAHBLTlOOI
=
CAHBLTOO1
;
else
CAHBLTlOOI
=
CAHBLTl10
;
end
CAHBLTOI1
:
begin
CAHBLTIOOI
=
"M2EXTEND"
;
CAHBLTO00
=
CAHBLTI11
;
if
(
CAHBLTII0
)
CAHBLTlOOI
=
CAHBLTII1
;
else
CAHBLTlOOI
=
CAHBLTOI1
;
end
CAHBLTIl1
:
begin
CAHBLTIOOI
=
"M3EXTEND"
;
CAHBLTO00
=
CAHBLTl11
;
if
(
CAHBLTII0
)
CAHBLTlOOI
=
CAHBLTll1
;
else
CAHBLTlOOI
=
CAHBLTIl1
;
end
CAHBLTO10
:
begin
CAHBLTIOOI
=
"M0LOCK"
;
if
(
CAHBLTlI0
)
if
(
CAHBLTOI0
[
0
]
)
begin
CAHBLTO00
=
CAHBLTl01
;
if
(
CAHBLTII0
)
CAHBLTlOOI
=
CAHBLTO10
;
else
CAHBLTlOOI
=
CAHBLTI10
;
end
else
CAHBLTlOOI
=
CAHBLTO10
;
else
CAHBLTlOOI
=
CAHBLTl00
;
end
CAHBLTI10
:
begin
CAHBLTIOOI
=
"M0LOCKEXTEND"
;
CAHBLTO00
=
CAHBLTl01
;
if
(
CAHBLTII0
)
CAHBLTlOOI
=
CAHBLTO10
;
else
CAHBLTlOOI
=
CAHBLTI10
;
end
CAHBLTIO1
:
begin
CAHBLTIOOI
=
"M1LOCK"
;
if
(
CAHBLTOl0
)
if
(
CAHBLTOI0
[
1
]
)
begin
CAHBLTO00
=
CAHBLTO11
;
if
(
CAHBLTII0
)
CAHBLTlOOI
=
CAHBLTIO1
;
else
CAHBLTlOOI
=
CAHBLTlO1
;
end
else
CAHBLTlOOI
=
CAHBLTIO1
;
else
CAHBLTlOOI
=
CAHBLTOO1
;
end
CAHBLTlO1
:
begin
CAHBLTIOOI
=
"M1LOCKEXTEND"
;
CAHBLTO00
=
CAHBLTO11
;
if
(
CAHBLTII0
)
CAHBLTlOOI
=
CAHBLTIO1
;
else
CAHBLTlOOI
=
CAHBLTlO1
;
end
CAHBLTlI1
:
begin
CAHBLTIOOI
=
"M2LOCK"
;
if
(
CAHBLTIl0
)
if
(
CAHBLTOI0
[
2
]
)
begin
CAHBLTO00
=
CAHBLTI11
;
if
(
CAHBLTII0
)
CAHBLTlOOI
=
CAHBLTlI1
;
else
CAHBLTlOOI
=
CAHBLTOl1
;
end
else
CAHBLTlOOI
=
CAHBLTlI1
;
else
CAHBLTlOOI
=
CAHBLTII1
;
end
CAHBLTOl1
:
begin
CAHBLTIOOI
=
"M2LOCKEXTEND"
;
CAHBLTO00
=
CAHBLTI11
;
if
(
CAHBLTII0
)
CAHBLTlOOI
=
CAHBLTlI1
;
else
CAHBLTlOOI
=
CAHBLTOl1
;
end
CAHBLTO01
:
begin
CAHBLTIOOI
=
"M3LOCK"
;
if
(
CAHBLTll0
)
if
(
CAHBLTOI0
[
3
]
)
begin
CAHBLTO00
=
CAHBLTl11
;
if
(
CAHBLTII0
)
CAHBLTlOOI
=
CAHBLTO01
;
else
CAHBLTlOOI
=
CAHBLTI01
;
end
else
CAHBLTlOOI
=
CAHBLTO01
;
else
CAHBLTlOOI
=
CAHBLTll1
;
end
CAHBLTI01
:
begin
CAHBLTIOOI
=
"M3LOCKEXTEND"
;
CAHBLTO00
=
CAHBLTl11
;
if
(
CAHBLTII0
)
CAHBLTlOOI
=
CAHBLTO01
;
else
CAHBLTlOOI
=
CAHBLTI01
;
end
default
:
CAHBLTlOOI
=
CAHBLTll1
;
endcase
end
always
@
(
posedge
HCLK
or
negedge
CAHBLTOO0
)
begin
if
(
(
!
CAHBLTOO0
)
||
(
!
CAHBLTIO0
)
)
CAHBLTOIOI
<=
CAHBLTll1
;
else
CAHBLTOIOI
<=
CAHBLTlOOI
;
end
endmodule
